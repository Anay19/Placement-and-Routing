magic
tech scmos
timestamp 11111111111
<< m1 >>
rect 73 5 74 6 
<< m2 >>
rect 73 5 74 6 
<< m2c >>
rect 73 5 74 6 
<< m1 >>
rect 73 5 74 6 
<< m2 >>
rect 73 5 74 6 
<< m1 >>
rect 74 5 75 6 
<< m1 >>
rect 75 5 76 6 
<< m1 >>
rect 76 5 77 6 
<< m1 >>
rect 77 5 78 6 
<< m1 >>
rect 78 5 79 6 
<< m1 >>
rect 79 5 80 6 
<< m1 >>
rect 80 5 81 6 
<< m1 >>
rect 81 5 82 6 
<< m1 >>
rect 82 5 83 6 
<< m1 >>
rect 83 5 84 6 
<< m1 >>
rect 84 5 85 6 
<< m1 >>
rect 85 5 86 6 
<< m1 >>
rect 86 5 87 6 
<< m1 >>
rect 87 5 88 6 
<< m1 >>
rect 88 5 89 6 
<< m1 >>
rect 89 5 90 6 
<< m1 >>
rect 90 5 91 6 
<< m1 >>
rect 91 5 92 6 
<< m1 >>
rect 92 5 93 6 
<< m1 >>
rect 93 5 94 6 
<< m1 >>
rect 94 5 95 6 
<< m1 >>
rect 95 5 96 6 
<< m1 >>
rect 96 5 97 6 
<< m1 >>
rect 97 5 98 6 
<< m1 >>
rect 98 5 99 6 
<< m1 >>
rect 99 5 100 6 
<< m1 >>
rect 100 5 101 6 
<< m1 >>
rect 101 5 102 6 
<< m1 >>
rect 102 5 103 6 
<< m1 >>
rect 103 5 104 6 
<< m1 >>
rect 104 5 105 6 
<< m1 >>
rect 105 5 106 6 
<< m1 >>
rect 106 5 107 6 
<< m1 >>
rect 107 5 108 6 
<< m1 >>
rect 108 5 109 6 
<< m1 >>
rect 109 5 110 6 
<< m1 >>
rect 110 5 111 6 
<< m1 >>
rect 111 5 112 6 
<< m1 >>
rect 112 5 113 6 
<< m1 >>
rect 113 5 114 6 
<< m1 >>
rect 114 5 115 6 
<< m1 >>
rect 115 5 116 6 
<< m1 >>
rect 116 5 117 6 
<< m1 >>
rect 117 5 118 6 
<< m1 >>
rect 118 5 119 6 
<< m1 >>
rect 119 5 120 6 
<< m1 >>
rect 120 5 121 6 
<< m1 >>
rect 121 5 122 6 
<< m1 >>
rect 122 5 123 6 
<< m1 >>
rect 123 5 124 6 
<< m1 >>
rect 124 5 125 6 
<< m1 >>
rect 125 5 126 6 
<< m1 >>
rect 126 5 127 6 
<< m1 >>
rect 127 5 128 6 
<< m1 >>
rect 128 5 129 6 
<< m2 >>
rect 128 5 129 6 
<< m2c >>
rect 128 5 129 6 
<< m1 >>
rect 128 5 129 6 
<< m2 >>
rect 128 5 129 6 
<< m2 >>
rect 73 6 74 7 
<< m2 >>
rect 128 6 129 7 
<< m1 >>
rect 37 7 38 8 
<< m2 >>
rect 37 7 38 8 
<< m1 >>
rect 38 7 39 8 
<< m2 >>
rect 38 7 39 8 
<< m1 >>
rect 39 7 40 8 
<< m2 >>
rect 39 7 40 8 
<< m1 >>
rect 40 7 41 8 
<< m2 >>
rect 40 7 41 8 
<< m1 >>
rect 41 7 42 8 
<< m2 >>
rect 41 7 42 8 
<< m1 >>
rect 42 7 43 8 
<< m2 >>
rect 42 7 43 8 
<< m1 >>
rect 43 7 44 8 
<< m2 >>
rect 43 7 44 8 
<< m1 >>
rect 44 7 45 8 
<< m2 >>
rect 44 7 45 8 
<< m1 >>
rect 45 7 46 8 
<< m2 >>
rect 45 7 46 8 
<< m1 >>
rect 46 7 47 8 
<< m2 >>
rect 46 7 47 8 
<< m1 >>
rect 47 7 48 8 
<< m2 >>
rect 47 7 48 8 
<< m1 >>
rect 48 7 49 8 
<< m2 >>
rect 48 7 49 8 
<< m1 >>
rect 49 7 50 8 
<< m2 >>
rect 49 7 50 8 
<< m1 >>
rect 50 7 51 8 
<< m2 >>
rect 50 7 51 8 
<< m1 >>
rect 51 7 52 8 
<< m1 >>
rect 52 7 53 8 
<< m1 >>
rect 53 7 54 8 
<< m1 >>
rect 54 7 55 8 
<< m1 >>
rect 55 7 56 8 
<< m1 >>
rect 56 7 57 8 
<< m1 >>
rect 57 7 58 8 
<< m1 >>
rect 58 7 59 8 
<< m1 >>
rect 59 7 60 8 
<< m1 >>
rect 60 7 61 8 
<< m1 >>
rect 61 7 62 8 
<< m1 >>
rect 62 7 63 8 
<< m1 >>
rect 63 7 64 8 
<< m1 >>
rect 64 7 65 8 
<< m1 >>
rect 65 7 66 8 
<< m1 >>
rect 66 7 67 8 
<< m1 >>
rect 67 7 68 8 
<< m1 >>
rect 68 7 69 8 
<< m1 >>
rect 69 7 70 8 
<< m1 >>
rect 70 7 71 8 
<< m1 >>
rect 71 7 72 8 
<< m1 >>
rect 72 7 73 8 
<< m1 >>
rect 73 7 74 8 
<< m2 >>
rect 73 7 74 8 
<< m1 >>
rect 74 7 75 8 
<< m1 >>
rect 75 7 76 8 
<< m1 >>
rect 76 7 77 8 
<< m1 >>
rect 77 7 78 8 
<< m1 >>
rect 78 7 79 8 
<< m1 >>
rect 79 7 80 8 
<< m1 >>
rect 80 7 81 8 
<< m1 >>
rect 81 7 82 8 
<< m1 >>
rect 82 7 83 8 
<< m1 >>
rect 83 7 84 8 
<< m1 >>
rect 84 7 85 8 
<< m1 >>
rect 85 7 86 8 
<< m1 >>
rect 86 7 87 8 
<< m1 >>
rect 87 7 88 8 
<< m1 >>
rect 88 7 89 8 
<< m1 >>
rect 89 7 90 8 
<< m1 >>
rect 90 7 91 8 
<< m1 >>
rect 91 7 92 8 
<< m2 >>
rect 91 7 92 8 
<< m1 >>
rect 92 7 93 8 
<< m2 >>
rect 92 7 93 8 
<< m1 >>
rect 93 7 94 8 
<< m2 >>
rect 93 7 94 8 
<< m1 >>
rect 94 7 95 8 
<< m2 >>
rect 94 7 95 8 
<< m1 >>
rect 95 7 96 8 
<< m2 >>
rect 95 7 96 8 
<< m1 >>
rect 96 7 97 8 
<< m2 >>
rect 96 7 97 8 
<< m1 >>
rect 97 7 98 8 
<< m2 >>
rect 97 7 98 8 
<< m1 >>
rect 98 7 99 8 
<< m2 >>
rect 98 7 99 8 
<< m1 >>
rect 99 7 100 8 
<< m2 >>
rect 99 7 100 8 
<< m1 >>
rect 100 7 101 8 
<< m2 >>
rect 100 7 101 8 
<< m1 >>
rect 101 7 102 8 
<< m2 >>
rect 101 7 102 8 
<< m1 >>
rect 102 7 103 8 
<< m2 >>
rect 102 7 103 8 
<< m1 >>
rect 103 7 104 8 
<< m2 >>
rect 103 7 104 8 
<< m1 >>
rect 104 7 105 8 
<< m2 >>
rect 104 7 105 8 
<< m1 >>
rect 105 7 106 8 
<< m2 >>
rect 105 7 106 8 
<< m1 >>
rect 106 7 107 8 
<< m2 >>
rect 106 7 107 8 
<< m1 >>
rect 107 7 108 8 
<< m2 >>
rect 107 7 108 8 
<< m1 >>
rect 108 7 109 8 
<< m2 >>
rect 108 7 109 8 
<< m1 >>
rect 109 7 110 8 
<< m2 >>
rect 109 7 110 8 
<< m1 >>
rect 110 7 111 8 
<< m2 >>
rect 110 7 111 8 
<< m1 >>
rect 111 7 112 8 
<< m2 >>
rect 111 7 112 8 
<< m1 >>
rect 112 7 113 8 
<< m2 >>
rect 112 7 113 8 
<< m1 >>
rect 113 7 114 8 
<< m2 >>
rect 113 7 114 8 
<< m1 >>
rect 114 7 115 8 
<< m2 >>
rect 114 7 115 8 
<< m1 >>
rect 115 7 116 8 
<< m2 >>
rect 115 7 116 8 
<< m1 >>
rect 116 7 117 8 
<< m2 >>
rect 116 7 117 8 
<< m1 >>
rect 117 7 118 8 
<< m2 >>
rect 117 7 118 8 
<< m1 >>
rect 118 7 119 8 
<< m2 >>
rect 118 7 119 8 
<< m1 >>
rect 119 7 120 8 
<< m2 >>
rect 119 7 120 8 
<< m1 >>
rect 120 7 121 8 
<< m2 >>
rect 120 7 121 8 
<< m1 >>
rect 121 7 122 8 
<< m2 >>
rect 121 7 122 8 
<< m1 >>
rect 122 7 123 8 
<< m2 >>
rect 122 7 123 8 
<< m1 >>
rect 123 7 124 8 
<< m2 >>
rect 123 7 124 8 
<< m1 >>
rect 124 7 125 8 
<< m2 >>
rect 124 7 125 8 
<< m2 >>
rect 125 7 126 8 
<< m1 >>
rect 126 7 127 8 
<< m2 >>
rect 126 7 127 8 
<< m2c >>
rect 126 7 127 8 
<< m1 >>
rect 126 7 127 8 
<< m2 >>
rect 126 7 127 8 
<< m1 >>
rect 127 7 128 8 
<< m1 >>
rect 128 7 129 8 
<< m2 >>
rect 128 7 129 8 
<< m1 >>
rect 129 7 130 8 
<< m1 >>
rect 130 7 131 8 
<< m1 >>
rect 131 7 132 8 
<< m1 >>
rect 132 7 133 8 
<< m1 >>
rect 133 7 134 8 
<< m1 >>
rect 134 7 135 8 
<< m1 >>
rect 135 7 136 8 
<< m1 >>
rect 136 7 137 8 
<< m1 >>
rect 137 7 138 8 
<< m1 >>
rect 138 7 139 8 
<< m1 >>
rect 139 7 140 8 
<< m1 >>
rect 140 7 141 8 
<< m1 >>
rect 141 7 142 8 
<< m1 >>
rect 142 7 143 8 
<< m1 >>
rect 37 8 38 9 
<< m2 >>
rect 37 8 38 9 
<< m2 >>
rect 50 8 51 9 
<< m2 >>
rect 73 8 74 9 
<< m2 >>
rect 91 8 92 9 
<< m1 >>
rect 124 8 125 9 
<< m2 >>
rect 128 8 129 9 
<< m1 >>
rect 142 8 143 9 
<< m1 >>
rect 37 9 38 10 
<< m2 >>
rect 37 9 38 10 
<< m1 >>
rect 50 9 51 10 
<< m2 >>
rect 50 9 51 10 
<< m2c >>
rect 50 9 51 10 
<< m1 >>
rect 50 9 51 10 
<< m2 >>
rect 50 9 51 10 
<< m1 >>
rect 51 9 52 10 
<< m1 >>
rect 52 9 53 10 
<< m1 >>
rect 73 9 74 10 
<< m2 >>
rect 73 9 74 10 
<< m2c >>
rect 73 9 74 10 
<< m1 >>
rect 73 9 74 10 
<< m2 >>
rect 73 9 74 10 
<< m1 >>
rect 91 9 92 10 
<< m2 >>
rect 91 9 92 10 
<< m2c >>
rect 91 9 92 10 
<< m1 >>
rect 91 9 92 10 
<< m2 >>
rect 91 9 92 10 
<< m1 >>
rect 124 9 125 10 
<< m1 >>
rect 128 9 129 10 
<< m2 >>
rect 128 9 129 10 
<< m2c >>
rect 128 9 129 10 
<< m1 >>
rect 128 9 129 10 
<< m2 >>
rect 128 9 129 10 
<< m1 >>
rect 142 9 143 10 
<< m1 >>
rect 37 10 38 11 
<< m2 >>
rect 37 10 38 11 
<< m1 >>
rect 52 10 53 11 
<< m1 >>
rect 73 10 74 11 
<< m1 >>
rect 91 10 92 11 
<< m1 >>
rect 124 10 125 11 
<< m1 >>
rect 128 10 129 11 
<< m1 >>
rect 142 10 143 11 
<< m1 >>
rect 37 11 38 12 
<< m2 >>
rect 37 11 38 12 
<< m1 >>
rect 52 11 53 12 
<< m1 >>
rect 73 11 74 12 
<< m1 >>
rect 91 11 92 12 
<< m1 >>
rect 124 11 125 12 
<< m1 >>
rect 128 11 129 12 
<< m1 >>
rect 142 11 143 12 
<< pdiffusion >>
rect 12 12 13 13 
<< pdiffusion >>
rect 13 12 14 13 
<< pdiffusion >>
rect 14 12 15 13 
<< pdiffusion >>
rect 15 12 16 13 
<< pdiffusion >>
rect 16 12 17 13 
<< pdiffusion >>
rect 17 12 18 13 
<< m1 >>
rect 37 12 38 13 
<< m2 >>
rect 37 12 38 13 
<< pdiffusion >>
rect 48 12 49 13 
<< pdiffusion >>
rect 49 12 50 13 
<< pdiffusion >>
rect 50 12 51 13 
<< pdiffusion >>
rect 51 12 52 13 
<< m1 >>
rect 52 12 53 13 
<< pdiffusion >>
rect 52 12 53 13 
<< pdiffusion >>
rect 53 12 54 13 
<< pdiffusion >>
rect 66 12 67 13 
<< pdiffusion >>
rect 67 12 68 13 
<< pdiffusion >>
rect 68 12 69 13 
<< pdiffusion >>
rect 69 12 70 13 
<< pdiffusion >>
rect 70 12 71 13 
<< pdiffusion >>
rect 71 12 72 13 
<< m1 >>
rect 73 12 74 13 
<< pdiffusion >>
rect 84 12 85 13 
<< pdiffusion >>
rect 85 12 86 13 
<< pdiffusion >>
rect 86 12 87 13 
<< pdiffusion >>
rect 87 12 88 13 
<< pdiffusion >>
rect 88 12 89 13 
<< pdiffusion >>
rect 89 12 90 13 
<< m1 >>
rect 91 12 92 13 
<< pdiffusion >>
rect 102 12 103 13 
<< pdiffusion >>
rect 103 12 104 13 
<< pdiffusion >>
rect 104 12 105 13 
<< pdiffusion >>
rect 105 12 106 13 
<< pdiffusion >>
rect 106 12 107 13 
<< pdiffusion >>
rect 107 12 108 13 
<< pdiffusion >>
rect 120 12 121 13 
<< pdiffusion >>
rect 121 12 122 13 
<< pdiffusion >>
rect 122 12 123 13 
<< pdiffusion >>
rect 123 12 124 13 
<< m1 >>
rect 124 12 125 13 
<< pdiffusion >>
rect 124 12 125 13 
<< pdiffusion >>
rect 125 12 126 13 
<< m1 >>
rect 128 12 129 13 
<< pdiffusion >>
rect 138 12 139 13 
<< pdiffusion >>
rect 139 12 140 13 
<< pdiffusion >>
rect 140 12 141 13 
<< pdiffusion >>
rect 141 12 142 13 
<< m1 >>
rect 142 12 143 13 
<< pdiffusion >>
rect 142 12 143 13 
<< pdiffusion >>
rect 143 12 144 13 
<< pdiffusion >>
rect 12 13 13 14 
<< pdiffusion >>
rect 13 13 14 14 
<< pdiffusion >>
rect 14 13 15 14 
<< pdiffusion >>
rect 15 13 16 14 
<< pdiffusion >>
rect 16 13 17 14 
<< pdiffusion >>
rect 17 13 18 14 
<< m1 >>
rect 37 13 38 14 
<< m2 >>
rect 37 13 38 14 
<< pdiffusion >>
rect 48 13 49 14 
<< pdiffusion >>
rect 49 13 50 14 
<< pdiffusion >>
rect 50 13 51 14 
<< pdiffusion >>
rect 51 13 52 14 
<< pdiffusion >>
rect 52 13 53 14 
<< pdiffusion >>
rect 53 13 54 14 
<< pdiffusion >>
rect 66 13 67 14 
<< pdiffusion >>
rect 67 13 68 14 
<< pdiffusion >>
rect 68 13 69 14 
<< pdiffusion >>
rect 69 13 70 14 
<< pdiffusion >>
rect 70 13 71 14 
<< pdiffusion >>
rect 71 13 72 14 
<< m1 >>
rect 73 13 74 14 
<< pdiffusion >>
rect 84 13 85 14 
<< pdiffusion >>
rect 85 13 86 14 
<< pdiffusion >>
rect 86 13 87 14 
<< pdiffusion >>
rect 87 13 88 14 
<< pdiffusion >>
rect 88 13 89 14 
<< pdiffusion >>
rect 89 13 90 14 
<< m1 >>
rect 91 13 92 14 
<< pdiffusion >>
rect 102 13 103 14 
<< pdiffusion >>
rect 103 13 104 14 
<< pdiffusion >>
rect 104 13 105 14 
<< pdiffusion >>
rect 105 13 106 14 
<< pdiffusion >>
rect 106 13 107 14 
<< pdiffusion >>
rect 107 13 108 14 
<< pdiffusion >>
rect 120 13 121 14 
<< pdiffusion >>
rect 121 13 122 14 
<< pdiffusion >>
rect 122 13 123 14 
<< pdiffusion >>
rect 123 13 124 14 
<< pdiffusion >>
rect 124 13 125 14 
<< pdiffusion >>
rect 125 13 126 14 
<< m1 >>
rect 128 13 129 14 
<< pdiffusion >>
rect 138 13 139 14 
<< pdiffusion >>
rect 139 13 140 14 
<< pdiffusion >>
rect 140 13 141 14 
<< pdiffusion >>
rect 141 13 142 14 
<< pdiffusion >>
rect 142 13 143 14 
<< pdiffusion >>
rect 143 13 144 14 
<< pdiffusion >>
rect 12 14 13 15 
<< pdiffusion >>
rect 13 14 14 15 
<< pdiffusion >>
rect 14 14 15 15 
<< pdiffusion >>
rect 15 14 16 15 
<< pdiffusion >>
rect 16 14 17 15 
<< pdiffusion >>
rect 17 14 18 15 
<< m1 >>
rect 37 14 38 15 
<< m2 >>
rect 37 14 38 15 
<< pdiffusion >>
rect 48 14 49 15 
<< pdiffusion >>
rect 49 14 50 15 
<< pdiffusion >>
rect 50 14 51 15 
<< pdiffusion >>
rect 51 14 52 15 
<< pdiffusion >>
rect 52 14 53 15 
<< pdiffusion >>
rect 53 14 54 15 
<< pdiffusion >>
rect 66 14 67 15 
<< pdiffusion >>
rect 67 14 68 15 
<< pdiffusion >>
rect 68 14 69 15 
<< pdiffusion >>
rect 69 14 70 15 
<< pdiffusion >>
rect 70 14 71 15 
<< pdiffusion >>
rect 71 14 72 15 
<< m1 >>
rect 73 14 74 15 
<< pdiffusion >>
rect 84 14 85 15 
<< pdiffusion >>
rect 85 14 86 15 
<< pdiffusion >>
rect 86 14 87 15 
<< pdiffusion >>
rect 87 14 88 15 
<< pdiffusion >>
rect 88 14 89 15 
<< pdiffusion >>
rect 89 14 90 15 
<< m1 >>
rect 91 14 92 15 
<< pdiffusion >>
rect 102 14 103 15 
<< pdiffusion >>
rect 103 14 104 15 
<< pdiffusion >>
rect 104 14 105 15 
<< pdiffusion >>
rect 105 14 106 15 
<< pdiffusion >>
rect 106 14 107 15 
<< pdiffusion >>
rect 107 14 108 15 
<< pdiffusion >>
rect 120 14 121 15 
<< pdiffusion >>
rect 121 14 122 15 
<< pdiffusion >>
rect 122 14 123 15 
<< pdiffusion >>
rect 123 14 124 15 
<< pdiffusion >>
rect 124 14 125 15 
<< pdiffusion >>
rect 125 14 126 15 
<< m1 >>
rect 128 14 129 15 
<< pdiffusion >>
rect 138 14 139 15 
<< pdiffusion >>
rect 139 14 140 15 
<< pdiffusion >>
rect 140 14 141 15 
<< pdiffusion >>
rect 141 14 142 15 
<< pdiffusion >>
rect 142 14 143 15 
<< pdiffusion >>
rect 143 14 144 15 
<< pdiffusion >>
rect 12 15 13 16 
<< pdiffusion >>
rect 13 15 14 16 
<< pdiffusion >>
rect 14 15 15 16 
<< pdiffusion >>
rect 15 15 16 16 
<< pdiffusion >>
rect 16 15 17 16 
<< pdiffusion >>
rect 17 15 18 16 
<< m1 >>
rect 37 15 38 16 
<< m2 >>
rect 37 15 38 16 
<< pdiffusion >>
rect 48 15 49 16 
<< pdiffusion >>
rect 49 15 50 16 
<< pdiffusion >>
rect 50 15 51 16 
<< pdiffusion >>
rect 51 15 52 16 
<< pdiffusion >>
rect 52 15 53 16 
<< pdiffusion >>
rect 53 15 54 16 
<< pdiffusion >>
rect 66 15 67 16 
<< pdiffusion >>
rect 67 15 68 16 
<< pdiffusion >>
rect 68 15 69 16 
<< pdiffusion >>
rect 69 15 70 16 
<< pdiffusion >>
rect 70 15 71 16 
<< pdiffusion >>
rect 71 15 72 16 
<< m1 >>
rect 73 15 74 16 
<< pdiffusion >>
rect 84 15 85 16 
<< pdiffusion >>
rect 85 15 86 16 
<< pdiffusion >>
rect 86 15 87 16 
<< pdiffusion >>
rect 87 15 88 16 
<< pdiffusion >>
rect 88 15 89 16 
<< pdiffusion >>
rect 89 15 90 16 
<< m1 >>
rect 91 15 92 16 
<< pdiffusion >>
rect 102 15 103 16 
<< pdiffusion >>
rect 103 15 104 16 
<< pdiffusion >>
rect 104 15 105 16 
<< pdiffusion >>
rect 105 15 106 16 
<< pdiffusion >>
rect 106 15 107 16 
<< pdiffusion >>
rect 107 15 108 16 
<< pdiffusion >>
rect 120 15 121 16 
<< pdiffusion >>
rect 121 15 122 16 
<< pdiffusion >>
rect 122 15 123 16 
<< pdiffusion >>
rect 123 15 124 16 
<< pdiffusion >>
rect 124 15 125 16 
<< pdiffusion >>
rect 125 15 126 16 
<< m1 >>
rect 128 15 129 16 
<< pdiffusion >>
rect 138 15 139 16 
<< pdiffusion >>
rect 139 15 140 16 
<< pdiffusion >>
rect 140 15 141 16 
<< pdiffusion >>
rect 141 15 142 16 
<< pdiffusion >>
rect 142 15 143 16 
<< pdiffusion >>
rect 143 15 144 16 
<< pdiffusion >>
rect 12 16 13 17 
<< pdiffusion >>
rect 13 16 14 17 
<< pdiffusion >>
rect 14 16 15 17 
<< pdiffusion >>
rect 15 16 16 17 
<< pdiffusion >>
rect 16 16 17 17 
<< pdiffusion >>
rect 17 16 18 17 
<< m1 >>
rect 37 16 38 17 
<< m2 >>
rect 37 16 38 17 
<< pdiffusion >>
rect 48 16 49 17 
<< pdiffusion >>
rect 49 16 50 17 
<< pdiffusion >>
rect 50 16 51 17 
<< pdiffusion >>
rect 51 16 52 17 
<< pdiffusion >>
rect 52 16 53 17 
<< pdiffusion >>
rect 53 16 54 17 
<< pdiffusion >>
rect 66 16 67 17 
<< pdiffusion >>
rect 67 16 68 17 
<< pdiffusion >>
rect 68 16 69 17 
<< pdiffusion >>
rect 69 16 70 17 
<< pdiffusion >>
rect 70 16 71 17 
<< pdiffusion >>
rect 71 16 72 17 
<< m1 >>
rect 73 16 74 17 
<< pdiffusion >>
rect 84 16 85 17 
<< pdiffusion >>
rect 85 16 86 17 
<< pdiffusion >>
rect 86 16 87 17 
<< pdiffusion >>
rect 87 16 88 17 
<< pdiffusion >>
rect 88 16 89 17 
<< pdiffusion >>
rect 89 16 90 17 
<< m1 >>
rect 91 16 92 17 
<< pdiffusion >>
rect 102 16 103 17 
<< pdiffusion >>
rect 103 16 104 17 
<< pdiffusion >>
rect 104 16 105 17 
<< pdiffusion >>
rect 105 16 106 17 
<< pdiffusion >>
rect 106 16 107 17 
<< pdiffusion >>
rect 107 16 108 17 
<< pdiffusion >>
rect 120 16 121 17 
<< pdiffusion >>
rect 121 16 122 17 
<< pdiffusion >>
rect 122 16 123 17 
<< pdiffusion >>
rect 123 16 124 17 
<< pdiffusion >>
rect 124 16 125 17 
<< pdiffusion >>
rect 125 16 126 17 
<< m1 >>
rect 128 16 129 17 
<< pdiffusion >>
rect 138 16 139 17 
<< pdiffusion >>
rect 139 16 140 17 
<< pdiffusion >>
rect 140 16 141 17 
<< pdiffusion >>
rect 141 16 142 17 
<< pdiffusion >>
rect 142 16 143 17 
<< pdiffusion >>
rect 143 16 144 17 
<< pdiffusion >>
rect 12 17 13 18 
<< pdiffusion >>
rect 13 17 14 18 
<< pdiffusion >>
rect 14 17 15 18 
<< pdiffusion >>
rect 15 17 16 18 
<< pdiffusion >>
rect 16 17 17 18 
<< pdiffusion >>
rect 17 17 18 18 
<< m1 >>
rect 37 17 38 18 
<< m2 >>
rect 37 17 38 18 
<< pdiffusion >>
rect 48 17 49 18 
<< m1 >>
rect 49 17 50 18 
<< pdiffusion >>
rect 49 17 50 18 
<< pdiffusion >>
rect 50 17 51 18 
<< pdiffusion >>
rect 51 17 52 18 
<< pdiffusion >>
rect 52 17 53 18 
<< pdiffusion >>
rect 53 17 54 18 
<< pdiffusion >>
rect 66 17 67 18 
<< m1 >>
rect 67 17 68 18 
<< pdiffusion >>
rect 67 17 68 18 
<< pdiffusion >>
rect 68 17 69 18 
<< pdiffusion >>
rect 69 17 70 18 
<< m1 >>
rect 70 17 71 18 
<< pdiffusion >>
rect 70 17 71 18 
<< pdiffusion >>
rect 71 17 72 18 
<< m1 >>
rect 73 17 74 18 
<< pdiffusion >>
rect 84 17 85 18 
<< pdiffusion >>
rect 85 17 86 18 
<< pdiffusion >>
rect 86 17 87 18 
<< pdiffusion >>
rect 87 17 88 18 
<< pdiffusion >>
rect 88 17 89 18 
<< pdiffusion >>
rect 89 17 90 18 
<< m1 >>
rect 91 17 92 18 
<< pdiffusion >>
rect 102 17 103 18 
<< m1 >>
rect 103 17 104 18 
<< pdiffusion >>
rect 103 17 104 18 
<< pdiffusion >>
rect 104 17 105 18 
<< pdiffusion >>
rect 105 17 106 18 
<< pdiffusion >>
rect 106 17 107 18 
<< pdiffusion >>
rect 107 17 108 18 
<< pdiffusion >>
rect 120 17 121 18 
<< pdiffusion >>
rect 121 17 122 18 
<< pdiffusion >>
rect 122 17 123 18 
<< pdiffusion >>
rect 123 17 124 18 
<< pdiffusion >>
rect 124 17 125 18 
<< pdiffusion >>
rect 125 17 126 18 
<< m1 >>
rect 128 17 129 18 
<< pdiffusion >>
rect 138 17 139 18 
<< pdiffusion >>
rect 139 17 140 18 
<< pdiffusion >>
rect 140 17 141 18 
<< pdiffusion >>
rect 141 17 142 18 
<< pdiffusion >>
rect 142 17 143 18 
<< pdiffusion >>
rect 143 17 144 18 
<< m1 >>
rect 37 18 38 19 
<< m2 >>
rect 37 18 38 19 
<< m1 >>
rect 49 18 50 19 
<< m1 >>
rect 67 18 68 19 
<< m1 >>
rect 70 18 71 19 
<< m1 >>
rect 73 18 74 19 
<< m1 >>
rect 91 18 92 19 
<< m1 >>
rect 103 18 104 19 
<< m1 >>
rect 128 18 129 19 
<< m1 >>
rect 37 19 38 20 
<< m2 >>
rect 37 19 38 20 
<< m1 >>
rect 49 19 50 20 
<< m1 >>
rect 67 19 68 20 
<< m1 >>
rect 70 19 71 20 
<< m1 >>
rect 73 19 74 20 
<< m1 >>
rect 91 19 92 20 
<< m1 >>
rect 103 19 104 20 
<< m1 >>
rect 128 19 129 20 
<< m1 >>
rect 37 20 38 21 
<< m2 >>
rect 37 20 38 21 
<< m1 >>
rect 49 20 50 21 
<< m1 >>
rect 50 20 51 21 
<< m1 >>
rect 51 20 52 21 
<< m1 >>
rect 52 20 53 21 
<< m1 >>
rect 53 20 54 21 
<< m1 >>
rect 54 20 55 21 
<< m1 >>
rect 55 20 56 21 
<< m1 >>
rect 56 20 57 21 
<< m1 >>
rect 57 20 58 21 
<< m1 >>
rect 58 20 59 21 
<< m1 >>
rect 59 20 60 21 
<< m1 >>
rect 60 20 61 21 
<< m1 >>
rect 61 20 62 21 
<< m1 >>
rect 62 20 63 21 
<< m1 >>
rect 63 20 64 21 
<< m1 >>
rect 64 20 65 21 
<< m1 >>
rect 65 20 66 21 
<< m1 >>
rect 66 20 67 21 
<< m1 >>
rect 67 20 68 21 
<< m1 >>
rect 70 20 71 21 
<< m1 >>
rect 73 20 74 21 
<< m2 >>
rect 73 20 74 21 
<< m2c >>
rect 73 20 74 21 
<< m1 >>
rect 73 20 74 21 
<< m2 >>
rect 73 20 74 21 
<< m1 >>
rect 91 20 92 21 
<< m2 >>
rect 91 20 92 21 
<< m2c >>
rect 91 20 92 21 
<< m1 >>
rect 91 20 92 21 
<< m2 >>
rect 91 20 92 21 
<< m1 >>
rect 103 20 104 21 
<< m1 >>
rect 128 20 129 21 
<< m1 >>
rect 37 21 38 22 
<< m2 >>
rect 37 21 38 22 
<< m1 >>
rect 70 21 71 22 
<< m2 >>
rect 73 21 74 22 
<< m2 >>
rect 91 21 92 22 
<< m1 >>
rect 103 21 104 22 
<< m1 >>
rect 128 21 129 22 
<< m1 >>
rect 37 22 38 23 
<< m2 >>
rect 37 22 38 23 
<< m1 >>
rect 70 22 71 23 
<< m1 >>
rect 71 22 72 23 
<< m1 >>
rect 72 22 73 23 
<< m1 >>
rect 73 22 74 23 
<< m2 >>
rect 73 22 74 23 
<< m1 >>
rect 74 22 75 23 
<< m1 >>
rect 75 22 76 23 
<< m1 >>
rect 76 22 77 23 
<< m1 >>
rect 77 22 78 23 
<< m1 >>
rect 78 22 79 23 
<< m1 >>
rect 79 22 80 23 
<< m1 >>
rect 80 22 81 23 
<< m1 >>
rect 81 22 82 23 
<< m1 >>
rect 82 22 83 23 
<< m1 >>
rect 83 22 84 23 
<< m1 >>
rect 84 22 85 23 
<< m1 >>
rect 85 22 86 23 
<< m1 >>
rect 86 22 87 23 
<< m1 >>
rect 87 22 88 23 
<< m1 >>
rect 88 22 89 23 
<< m1 >>
rect 89 22 90 23 
<< m1 >>
rect 90 22 91 23 
<< m1 >>
rect 91 22 92 23 
<< m2 >>
rect 91 22 92 23 
<< m1 >>
rect 92 22 93 23 
<< m1 >>
rect 93 22 94 23 
<< m1 >>
rect 94 22 95 23 
<< m1 >>
rect 95 22 96 23 
<< m1 >>
rect 96 22 97 23 
<< m1 >>
rect 97 22 98 23 
<< m1 >>
rect 98 22 99 23 
<< m1 >>
rect 99 22 100 23 
<< m1 >>
rect 100 22 101 23 
<< m1 >>
rect 101 22 102 23 
<< m1 >>
rect 102 22 103 23 
<< m1 >>
rect 103 22 104 23 
<< m1 >>
rect 128 22 129 23 
<< m1 >>
rect 37 23 38 24 
<< m2 >>
rect 37 23 38 24 
<< m2 >>
rect 73 23 74 24 
<< m2 >>
rect 91 23 92 24 
<< m1 >>
rect 128 23 129 24 
<< m1 >>
rect 37 24 38 25 
<< m2 >>
rect 37 24 38 25 
<< m2 >>
rect 73 24 74 25 
<< m2 >>
rect 91 24 92 25 
<< m1 >>
rect 128 24 129 25 
<< m1 >>
rect 37 25 38 26 
<< m2 >>
rect 37 25 38 26 
<< m1 >>
rect 55 25 56 26 
<< m1 >>
rect 56 25 57 26 
<< m1 >>
rect 57 25 58 26 
<< m1 >>
rect 58 25 59 26 
<< m1 >>
rect 59 25 60 26 
<< m1 >>
rect 60 25 61 26 
<< m1 >>
rect 61 25 62 26 
<< m1 >>
rect 62 25 63 26 
<< m1 >>
rect 63 25 64 26 
<< m1 >>
rect 64 25 65 26 
<< m1 >>
rect 65 25 66 26 
<< m1 >>
rect 66 25 67 26 
<< m2 >>
rect 66 25 67 26 
<< m1 >>
rect 67 25 68 26 
<< m2 >>
rect 67 25 68 26 
<< m1 >>
rect 68 25 69 26 
<< m2 >>
rect 68 25 69 26 
<< m1 >>
rect 69 25 70 26 
<< m2 >>
rect 69 25 70 26 
<< m1 >>
rect 70 25 71 26 
<< m2 >>
rect 70 25 71 26 
<< m1 >>
rect 71 25 72 26 
<< m1 >>
rect 72 25 73 26 
<< m1 >>
rect 73 25 74 26 
<< m2 >>
rect 73 25 74 26 
<< m1 >>
rect 74 25 75 26 
<< m1 >>
rect 75 25 76 26 
<< m1 >>
rect 76 25 77 26 
<< m1 >>
rect 77 25 78 26 
<< m1 >>
rect 78 25 79 26 
<< m1 >>
rect 79 25 80 26 
<< m1 >>
rect 80 25 81 26 
<< m1 >>
rect 81 25 82 26 
<< m1 >>
rect 82 25 83 26 
<< m1 >>
rect 83 25 84 26 
<< m1 >>
rect 84 25 85 26 
<< m1 >>
rect 85 25 86 26 
<< m1 >>
rect 88 25 89 26 
<< m1 >>
rect 89 25 90 26 
<< m1 >>
rect 90 25 91 26 
<< m1 >>
rect 91 25 92 26 
<< m2 >>
rect 91 25 92 26 
<< m1 >>
rect 92 25 93 26 
<< m1 >>
rect 93 25 94 26 
<< m1 >>
rect 94 25 95 26 
<< m1 >>
rect 95 25 96 26 
<< m1 >>
rect 96 25 97 26 
<< m1 >>
rect 97 25 98 26 
<< m1 >>
rect 98 25 99 26 
<< m1 >>
rect 99 25 100 26 
<< m1 >>
rect 100 25 101 26 
<< m1 >>
rect 101 25 102 26 
<< m1 >>
rect 102 25 103 26 
<< m1 >>
rect 103 25 104 26 
<< m1 >>
rect 104 25 105 26 
<< m1 >>
rect 105 25 106 26 
<< m1 >>
rect 106 25 107 26 
<< m1 >>
rect 107 25 108 26 
<< m1 >>
rect 108 25 109 26 
<< m1 >>
rect 109 25 110 26 
<< m1 >>
rect 110 25 111 26 
<< m1 >>
rect 111 25 112 26 
<< m1 >>
rect 112 25 113 26 
<< m1 >>
rect 113 25 114 26 
<< m1 >>
rect 114 25 115 26 
<< m1 >>
rect 115 25 116 26 
<< m1 >>
rect 116 25 117 26 
<< m1 >>
rect 117 25 118 26 
<< m1 >>
rect 118 25 119 26 
<< m1 >>
rect 119 25 120 26 
<< m1 >>
rect 120 25 121 26 
<< m1 >>
rect 121 25 122 26 
<< m1 >>
rect 122 25 123 26 
<< m1 >>
rect 123 25 124 26 
<< m1 >>
rect 124 25 125 26 
<< m1 >>
rect 128 25 129 26 
<< m1 >>
rect 37 26 38 27 
<< m2 >>
rect 37 26 38 27 
<< m1 >>
rect 55 26 56 27 
<< m2 >>
rect 66 26 67 27 
<< m2 >>
rect 70 26 71 27 
<< m2 >>
rect 73 26 74 27 
<< m1 >>
rect 85 26 86 27 
<< m1 >>
rect 88 26 89 27 
<< m2 >>
rect 91 26 92 27 
<< m1 >>
rect 124 26 125 27 
<< m1 >>
rect 128 26 129 27 
<< m1 >>
rect 13 27 14 28 
<< m1 >>
rect 14 27 15 28 
<< m1 >>
rect 15 27 16 28 
<< m1 >>
rect 16 27 17 28 
<< m1 >>
rect 17 27 18 28 
<< m1 >>
rect 18 27 19 28 
<< m1 >>
rect 19 27 20 28 
<< m1 >>
rect 37 27 38 28 
<< m2 >>
rect 37 27 38 28 
<< m1 >>
rect 55 27 56 28 
<< m1 >>
rect 64 27 65 28 
<< m1 >>
rect 65 27 66 28 
<< m1 >>
rect 66 27 67 28 
<< m2 >>
rect 66 27 67 28 
<< m2c >>
rect 66 27 67 28 
<< m1 >>
rect 66 27 67 28 
<< m2 >>
rect 66 27 67 28 
<< m1 >>
rect 70 27 71 28 
<< m2 >>
rect 70 27 71 28 
<< m2c >>
rect 70 27 71 28 
<< m1 >>
rect 70 27 71 28 
<< m2 >>
rect 70 27 71 28 
<< m1 >>
rect 73 27 74 28 
<< m2 >>
rect 73 27 74 28 
<< m2c >>
rect 73 27 74 28 
<< m1 >>
rect 73 27 74 28 
<< m2 >>
rect 73 27 74 28 
<< m1 >>
rect 85 27 86 28 
<< m1 >>
rect 88 27 89 28 
<< m1 >>
rect 91 27 92 28 
<< m2 >>
rect 91 27 92 28 
<< m2c >>
rect 91 27 92 28 
<< m1 >>
rect 91 27 92 28 
<< m2 >>
rect 91 27 92 28 
<< m1 >>
rect 124 27 125 28 
<< m1 >>
rect 128 27 129 28 
<< m1 >>
rect 13 28 14 29 
<< m2 >>
rect 16 28 17 29 
<< m2 >>
rect 17 28 18 29 
<< m2 >>
rect 18 28 19 29 
<< m1 >>
rect 19 28 20 29 
<< m2 >>
rect 19 28 20 29 
<< m1 >>
rect 37 28 38 29 
<< m2 >>
rect 37 28 38 29 
<< m1 >>
rect 52 28 53 29 
<< m1 >>
rect 53 28 54 29 
<< m2 >>
rect 53 28 54 29 
<< m2c >>
rect 53 28 54 29 
<< m1 >>
rect 53 28 54 29 
<< m2 >>
rect 53 28 54 29 
<< m2 >>
rect 54 28 55 29 
<< m1 >>
rect 55 28 56 29 
<< m2 >>
rect 55 28 56 29 
<< m1 >>
rect 64 28 65 29 
<< m1 >>
rect 70 28 71 29 
<< m1 >>
rect 73 28 74 29 
<< m1 >>
rect 85 28 86 29 
<< m1 >>
rect 88 28 89 29 
<< m1 >>
rect 91 28 92 29 
<< m1 >>
rect 124 28 125 29 
<< m1 >>
rect 128 28 129 29 
<< m1 >>
rect 13 29 14 30 
<< m1 >>
rect 16 29 17 30 
<< m2 >>
rect 16 29 17 30 
<< m1 >>
rect 19 29 20 30 
<< m2 >>
rect 19 29 20 30 
<< m1 >>
rect 37 29 38 30 
<< m2 >>
rect 37 29 38 30 
<< m1 >>
rect 52 29 53 30 
<< m1 >>
rect 55 29 56 30 
<< m2 >>
rect 55 29 56 30 
<< m1 >>
rect 64 29 65 30 
<< m1 >>
rect 70 29 71 30 
<< m1 >>
rect 73 29 74 30 
<< m1 >>
rect 85 29 86 30 
<< m1 >>
rect 88 29 89 30 
<< m1 >>
rect 91 29 92 30 
<< m1 >>
rect 124 29 125 30 
<< m1 >>
rect 128 29 129 30 
<< pdiffusion >>
rect 12 30 13 31 
<< m1 >>
rect 13 30 14 31 
<< pdiffusion >>
rect 13 30 14 31 
<< pdiffusion >>
rect 14 30 15 31 
<< m1 >>
rect 15 30 16 31 
<< m2 >>
rect 15 30 16 31 
<< m2c >>
rect 15 30 16 31 
<< m1 >>
rect 15 30 16 31 
<< m2 >>
rect 15 30 16 31 
<< pdiffusion >>
rect 15 30 16 31 
<< m1 >>
rect 16 30 17 31 
<< pdiffusion >>
rect 16 30 17 31 
<< pdiffusion >>
rect 17 30 18 31 
<< m1 >>
rect 19 30 20 31 
<< m2 >>
rect 19 30 20 31 
<< pdiffusion >>
rect 30 30 31 31 
<< pdiffusion >>
rect 31 30 32 31 
<< pdiffusion >>
rect 32 30 33 31 
<< pdiffusion >>
rect 33 30 34 31 
<< pdiffusion >>
rect 34 30 35 31 
<< pdiffusion >>
rect 35 30 36 31 
<< m1 >>
rect 37 30 38 31 
<< m2 >>
rect 37 30 38 31 
<< pdiffusion >>
rect 48 30 49 31 
<< pdiffusion >>
rect 49 30 50 31 
<< pdiffusion >>
rect 50 30 51 31 
<< pdiffusion >>
rect 51 30 52 31 
<< m1 >>
rect 52 30 53 31 
<< pdiffusion >>
rect 52 30 53 31 
<< pdiffusion >>
rect 53 30 54 31 
<< m1 >>
rect 55 30 56 31 
<< m2 >>
rect 55 30 56 31 
<< m1 >>
rect 64 30 65 31 
<< pdiffusion >>
rect 66 30 67 31 
<< pdiffusion >>
rect 67 30 68 31 
<< pdiffusion >>
rect 68 30 69 31 
<< pdiffusion >>
rect 69 30 70 31 
<< m1 >>
rect 70 30 71 31 
<< pdiffusion >>
rect 70 30 71 31 
<< pdiffusion >>
rect 71 30 72 31 
<< m1 >>
rect 73 30 74 31 
<< pdiffusion >>
rect 84 30 85 31 
<< m1 >>
rect 85 30 86 31 
<< pdiffusion >>
rect 85 30 86 31 
<< pdiffusion >>
rect 86 30 87 31 
<< pdiffusion >>
rect 87 30 88 31 
<< m1 >>
rect 88 30 89 31 
<< pdiffusion >>
rect 88 30 89 31 
<< pdiffusion >>
rect 89 30 90 31 
<< m1 >>
rect 91 30 92 31 
<< pdiffusion >>
rect 102 30 103 31 
<< pdiffusion >>
rect 103 30 104 31 
<< pdiffusion >>
rect 104 30 105 31 
<< pdiffusion >>
rect 105 30 106 31 
<< pdiffusion >>
rect 106 30 107 31 
<< pdiffusion >>
rect 107 30 108 31 
<< pdiffusion >>
rect 120 30 121 31 
<< pdiffusion >>
rect 121 30 122 31 
<< pdiffusion >>
rect 122 30 123 31 
<< pdiffusion >>
rect 123 30 124 31 
<< m1 >>
rect 124 30 125 31 
<< pdiffusion >>
rect 124 30 125 31 
<< pdiffusion >>
rect 125 30 126 31 
<< m1 >>
rect 128 30 129 31 
<< pdiffusion >>
rect 12 31 13 32 
<< pdiffusion >>
rect 13 31 14 32 
<< pdiffusion >>
rect 14 31 15 32 
<< pdiffusion >>
rect 15 31 16 32 
<< pdiffusion >>
rect 16 31 17 32 
<< pdiffusion >>
rect 17 31 18 32 
<< m1 >>
rect 19 31 20 32 
<< m2 >>
rect 19 31 20 32 
<< pdiffusion >>
rect 30 31 31 32 
<< pdiffusion >>
rect 31 31 32 32 
<< pdiffusion >>
rect 32 31 33 32 
<< pdiffusion >>
rect 33 31 34 32 
<< pdiffusion >>
rect 34 31 35 32 
<< pdiffusion >>
rect 35 31 36 32 
<< m1 >>
rect 37 31 38 32 
<< m2 >>
rect 37 31 38 32 
<< pdiffusion >>
rect 48 31 49 32 
<< pdiffusion >>
rect 49 31 50 32 
<< pdiffusion >>
rect 50 31 51 32 
<< pdiffusion >>
rect 51 31 52 32 
<< pdiffusion >>
rect 52 31 53 32 
<< pdiffusion >>
rect 53 31 54 32 
<< m1 >>
rect 55 31 56 32 
<< m2 >>
rect 55 31 56 32 
<< m1 >>
rect 64 31 65 32 
<< pdiffusion >>
rect 66 31 67 32 
<< pdiffusion >>
rect 67 31 68 32 
<< pdiffusion >>
rect 68 31 69 32 
<< pdiffusion >>
rect 69 31 70 32 
<< pdiffusion >>
rect 70 31 71 32 
<< pdiffusion >>
rect 71 31 72 32 
<< m1 >>
rect 73 31 74 32 
<< pdiffusion >>
rect 84 31 85 32 
<< pdiffusion >>
rect 85 31 86 32 
<< pdiffusion >>
rect 86 31 87 32 
<< pdiffusion >>
rect 87 31 88 32 
<< pdiffusion >>
rect 88 31 89 32 
<< pdiffusion >>
rect 89 31 90 32 
<< m1 >>
rect 91 31 92 32 
<< pdiffusion >>
rect 102 31 103 32 
<< pdiffusion >>
rect 103 31 104 32 
<< pdiffusion >>
rect 104 31 105 32 
<< pdiffusion >>
rect 105 31 106 32 
<< pdiffusion >>
rect 106 31 107 32 
<< pdiffusion >>
rect 107 31 108 32 
<< pdiffusion >>
rect 120 31 121 32 
<< pdiffusion >>
rect 121 31 122 32 
<< pdiffusion >>
rect 122 31 123 32 
<< pdiffusion >>
rect 123 31 124 32 
<< pdiffusion >>
rect 124 31 125 32 
<< pdiffusion >>
rect 125 31 126 32 
<< m1 >>
rect 128 31 129 32 
<< pdiffusion >>
rect 12 32 13 33 
<< pdiffusion >>
rect 13 32 14 33 
<< pdiffusion >>
rect 14 32 15 33 
<< pdiffusion >>
rect 15 32 16 33 
<< pdiffusion >>
rect 16 32 17 33 
<< pdiffusion >>
rect 17 32 18 33 
<< m1 >>
rect 19 32 20 33 
<< m2 >>
rect 19 32 20 33 
<< pdiffusion >>
rect 30 32 31 33 
<< pdiffusion >>
rect 31 32 32 33 
<< pdiffusion >>
rect 32 32 33 33 
<< pdiffusion >>
rect 33 32 34 33 
<< pdiffusion >>
rect 34 32 35 33 
<< pdiffusion >>
rect 35 32 36 33 
<< m1 >>
rect 37 32 38 33 
<< m2 >>
rect 37 32 38 33 
<< pdiffusion >>
rect 48 32 49 33 
<< pdiffusion >>
rect 49 32 50 33 
<< pdiffusion >>
rect 50 32 51 33 
<< pdiffusion >>
rect 51 32 52 33 
<< pdiffusion >>
rect 52 32 53 33 
<< pdiffusion >>
rect 53 32 54 33 
<< m1 >>
rect 55 32 56 33 
<< m2 >>
rect 55 32 56 33 
<< m1 >>
rect 64 32 65 33 
<< pdiffusion >>
rect 66 32 67 33 
<< pdiffusion >>
rect 67 32 68 33 
<< pdiffusion >>
rect 68 32 69 33 
<< pdiffusion >>
rect 69 32 70 33 
<< pdiffusion >>
rect 70 32 71 33 
<< pdiffusion >>
rect 71 32 72 33 
<< m1 >>
rect 73 32 74 33 
<< pdiffusion >>
rect 84 32 85 33 
<< pdiffusion >>
rect 85 32 86 33 
<< pdiffusion >>
rect 86 32 87 33 
<< pdiffusion >>
rect 87 32 88 33 
<< pdiffusion >>
rect 88 32 89 33 
<< pdiffusion >>
rect 89 32 90 33 
<< m1 >>
rect 91 32 92 33 
<< pdiffusion >>
rect 102 32 103 33 
<< pdiffusion >>
rect 103 32 104 33 
<< pdiffusion >>
rect 104 32 105 33 
<< pdiffusion >>
rect 105 32 106 33 
<< pdiffusion >>
rect 106 32 107 33 
<< pdiffusion >>
rect 107 32 108 33 
<< pdiffusion >>
rect 120 32 121 33 
<< pdiffusion >>
rect 121 32 122 33 
<< pdiffusion >>
rect 122 32 123 33 
<< pdiffusion >>
rect 123 32 124 33 
<< pdiffusion >>
rect 124 32 125 33 
<< pdiffusion >>
rect 125 32 126 33 
<< m1 >>
rect 128 32 129 33 
<< pdiffusion >>
rect 12 33 13 34 
<< pdiffusion >>
rect 13 33 14 34 
<< pdiffusion >>
rect 14 33 15 34 
<< pdiffusion >>
rect 15 33 16 34 
<< pdiffusion >>
rect 16 33 17 34 
<< pdiffusion >>
rect 17 33 18 34 
<< m1 >>
rect 19 33 20 34 
<< m2 >>
rect 19 33 20 34 
<< pdiffusion >>
rect 30 33 31 34 
<< pdiffusion >>
rect 31 33 32 34 
<< pdiffusion >>
rect 32 33 33 34 
<< pdiffusion >>
rect 33 33 34 34 
<< pdiffusion >>
rect 34 33 35 34 
<< pdiffusion >>
rect 35 33 36 34 
<< m1 >>
rect 37 33 38 34 
<< m2 >>
rect 37 33 38 34 
<< pdiffusion >>
rect 48 33 49 34 
<< pdiffusion >>
rect 49 33 50 34 
<< pdiffusion >>
rect 50 33 51 34 
<< pdiffusion >>
rect 51 33 52 34 
<< pdiffusion >>
rect 52 33 53 34 
<< pdiffusion >>
rect 53 33 54 34 
<< m1 >>
rect 55 33 56 34 
<< m2 >>
rect 55 33 56 34 
<< m1 >>
rect 64 33 65 34 
<< pdiffusion >>
rect 66 33 67 34 
<< pdiffusion >>
rect 67 33 68 34 
<< pdiffusion >>
rect 68 33 69 34 
<< pdiffusion >>
rect 69 33 70 34 
<< pdiffusion >>
rect 70 33 71 34 
<< pdiffusion >>
rect 71 33 72 34 
<< m1 >>
rect 73 33 74 34 
<< pdiffusion >>
rect 84 33 85 34 
<< pdiffusion >>
rect 85 33 86 34 
<< pdiffusion >>
rect 86 33 87 34 
<< pdiffusion >>
rect 87 33 88 34 
<< pdiffusion >>
rect 88 33 89 34 
<< pdiffusion >>
rect 89 33 90 34 
<< m1 >>
rect 91 33 92 34 
<< pdiffusion >>
rect 102 33 103 34 
<< pdiffusion >>
rect 103 33 104 34 
<< pdiffusion >>
rect 104 33 105 34 
<< pdiffusion >>
rect 105 33 106 34 
<< pdiffusion >>
rect 106 33 107 34 
<< pdiffusion >>
rect 107 33 108 34 
<< pdiffusion >>
rect 120 33 121 34 
<< pdiffusion >>
rect 121 33 122 34 
<< pdiffusion >>
rect 122 33 123 34 
<< pdiffusion >>
rect 123 33 124 34 
<< pdiffusion >>
rect 124 33 125 34 
<< pdiffusion >>
rect 125 33 126 34 
<< m1 >>
rect 128 33 129 34 
<< pdiffusion >>
rect 12 34 13 35 
<< pdiffusion >>
rect 13 34 14 35 
<< pdiffusion >>
rect 14 34 15 35 
<< pdiffusion >>
rect 15 34 16 35 
<< pdiffusion >>
rect 16 34 17 35 
<< pdiffusion >>
rect 17 34 18 35 
<< m1 >>
rect 19 34 20 35 
<< m2 >>
rect 19 34 20 35 
<< pdiffusion >>
rect 30 34 31 35 
<< pdiffusion >>
rect 31 34 32 35 
<< pdiffusion >>
rect 32 34 33 35 
<< pdiffusion >>
rect 33 34 34 35 
<< pdiffusion >>
rect 34 34 35 35 
<< pdiffusion >>
rect 35 34 36 35 
<< m1 >>
rect 37 34 38 35 
<< m2 >>
rect 37 34 38 35 
<< pdiffusion >>
rect 48 34 49 35 
<< pdiffusion >>
rect 49 34 50 35 
<< pdiffusion >>
rect 50 34 51 35 
<< pdiffusion >>
rect 51 34 52 35 
<< pdiffusion >>
rect 52 34 53 35 
<< pdiffusion >>
rect 53 34 54 35 
<< m1 >>
rect 55 34 56 35 
<< m2 >>
rect 55 34 56 35 
<< m1 >>
rect 64 34 65 35 
<< pdiffusion >>
rect 66 34 67 35 
<< pdiffusion >>
rect 67 34 68 35 
<< pdiffusion >>
rect 68 34 69 35 
<< pdiffusion >>
rect 69 34 70 35 
<< pdiffusion >>
rect 70 34 71 35 
<< pdiffusion >>
rect 71 34 72 35 
<< m1 >>
rect 73 34 74 35 
<< pdiffusion >>
rect 84 34 85 35 
<< pdiffusion >>
rect 85 34 86 35 
<< pdiffusion >>
rect 86 34 87 35 
<< pdiffusion >>
rect 87 34 88 35 
<< pdiffusion >>
rect 88 34 89 35 
<< pdiffusion >>
rect 89 34 90 35 
<< m1 >>
rect 91 34 92 35 
<< pdiffusion >>
rect 102 34 103 35 
<< pdiffusion >>
rect 103 34 104 35 
<< pdiffusion >>
rect 104 34 105 35 
<< pdiffusion >>
rect 105 34 106 35 
<< pdiffusion >>
rect 106 34 107 35 
<< pdiffusion >>
rect 107 34 108 35 
<< pdiffusion >>
rect 120 34 121 35 
<< pdiffusion >>
rect 121 34 122 35 
<< pdiffusion >>
rect 122 34 123 35 
<< pdiffusion >>
rect 123 34 124 35 
<< pdiffusion >>
rect 124 34 125 35 
<< pdiffusion >>
rect 125 34 126 35 
<< m1 >>
rect 128 34 129 35 
<< pdiffusion >>
rect 12 35 13 36 
<< m1 >>
rect 13 35 14 36 
<< pdiffusion >>
rect 13 35 14 36 
<< pdiffusion >>
rect 14 35 15 36 
<< pdiffusion >>
rect 15 35 16 36 
<< pdiffusion >>
rect 16 35 17 36 
<< pdiffusion >>
rect 17 35 18 36 
<< m1 >>
rect 19 35 20 36 
<< m2 >>
rect 19 35 20 36 
<< pdiffusion >>
rect 30 35 31 36 
<< m1 >>
rect 31 35 32 36 
<< pdiffusion >>
rect 31 35 32 36 
<< pdiffusion >>
rect 32 35 33 36 
<< m1 >>
rect 33 35 34 36 
<< m2 >>
rect 33 35 34 36 
<< m2c >>
rect 33 35 34 36 
<< m1 >>
rect 33 35 34 36 
<< m2 >>
rect 33 35 34 36 
<< pdiffusion >>
rect 33 35 34 36 
<< m1 >>
rect 34 35 35 36 
<< pdiffusion >>
rect 34 35 35 36 
<< pdiffusion >>
rect 35 35 36 36 
<< m1 >>
rect 37 35 38 36 
<< m2 >>
rect 37 35 38 36 
<< pdiffusion >>
rect 48 35 49 36 
<< pdiffusion >>
rect 49 35 50 36 
<< pdiffusion >>
rect 50 35 51 36 
<< pdiffusion >>
rect 51 35 52 36 
<< m1 >>
rect 52 35 53 36 
<< pdiffusion >>
rect 52 35 53 36 
<< pdiffusion >>
rect 53 35 54 36 
<< m1 >>
rect 55 35 56 36 
<< m2 >>
rect 55 35 56 36 
<< m1 >>
rect 64 35 65 36 
<< pdiffusion >>
rect 66 35 67 36 
<< pdiffusion >>
rect 67 35 68 36 
<< pdiffusion >>
rect 68 35 69 36 
<< pdiffusion >>
rect 69 35 70 36 
<< pdiffusion >>
rect 70 35 71 36 
<< pdiffusion >>
rect 71 35 72 36 
<< m1 >>
rect 73 35 74 36 
<< pdiffusion >>
rect 84 35 85 36 
<< pdiffusion >>
rect 85 35 86 36 
<< pdiffusion >>
rect 86 35 87 36 
<< pdiffusion >>
rect 87 35 88 36 
<< pdiffusion >>
rect 88 35 89 36 
<< pdiffusion >>
rect 89 35 90 36 
<< m1 >>
rect 91 35 92 36 
<< pdiffusion >>
rect 102 35 103 36 
<< m1 >>
rect 103 35 104 36 
<< pdiffusion >>
rect 103 35 104 36 
<< pdiffusion >>
rect 104 35 105 36 
<< pdiffusion >>
rect 105 35 106 36 
<< pdiffusion >>
rect 106 35 107 36 
<< pdiffusion >>
rect 107 35 108 36 
<< pdiffusion >>
rect 120 35 121 36 
<< m1 >>
rect 121 35 122 36 
<< pdiffusion >>
rect 121 35 122 36 
<< pdiffusion >>
rect 122 35 123 36 
<< pdiffusion >>
rect 123 35 124 36 
<< pdiffusion >>
rect 124 35 125 36 
<< pdiffusion >>
rect 125 35 126 36 
<< m1 >>
rect 128 35 129 36 
<< m1 >>
rect 13 36 14 37 
<< m1 >>
rect 19 36 20 37 
<< m2 >>
rect 19 36 20 37 
<< m1 >>
rect 31 36 32 37 
<< m1 >>
rect 34 36 35 37 
<< m2 >>
rect 34 36 35 37 
<< m1 >>
rect 37 36 38 37 
<< m2 >>
rect 37 36 38 37 
<< m1 >>
rect 52 36 53 37 
<< m1 >>
rect 55 36 56 37 
<< m2 >>
rect 55 36 56 37 
<< m1 >>
rect 64 36 65 37 
<< m1 >>
rect 73 36 74 37 
<< m1 >>
rect 91 36 92 37 
<< m1 >>
rect 103 36 104 37 
<< m1 >>
rect 121 36 122 37 
<< m1 >>
rect 128 36 129 37 
<< m1 >>
rect 13 37 14 38 
<< m1 >>
rect 19 37 20 38 
<< m2 >>
rect 19 37 20 38 
<< m1 >>
rect 31 37 32 38 
<< m2 >>
rect 34 37 35 38 
<< m2 >>
rect 35 37 36 38 
<< m2 >>
rect 36 37 37 38 
<< m1 >>
rect 37 37 38 38 
<< m2 >>
rect 37 37 38 38 
<< m1 >>
rect 52 37 53 38 
<< m1 >>
rect 53 37 54 38 
<< m1 >>
rect 54 37 55 38 
<< m1 >>
rect 55 37 56 38 
<< m2 >>
rect 55 37 56 38 
<< m1 >>
rect 64 37 65 38 
<< m1 >>
rect 73 37 74 38 
<< m1 >>
rect 91 37 92 38 
<< m1 >>
rect 100 37 101 38 
<< m1 >>
rect 101 37 102 38 
<< m1 >>
rect 102 37 103 38 
<< m1 >>
rect 103 37 104 38 
<< m1 >>
rect 121 37 122 38 
<< m1 >>
rect 128 37 129 38 
<< m1 >>
rect 13 38 14 39 
<< m1 >>
rect 19 38 20 39 
<< m2 >>
rect 19 38 20 39 
<< m1 >>
rect 31 38 32 39 
<< m1 >>
rect 32 38 33 39 
<< m1 >>
rect 33 38 34 39 
<< m1 >>
rect 34 38 35 39 
<< m1 >>
rect 35 38 36 39 
<< m1 >>
rect 36 38 37 39 
<< m1 >>
rect 37 38 38 39 
<< m2 >>
rect 55 38 56 39 
<< m1 >>
rect 64 38 65 39 
<< m1 >>
rect 73 38 74 39 
<< m1 >>
rect 91 38 92 39 
<< m1 >>
rect 100 38 101 39 
<< m1 >>
rect 121 38 122 39 
<< m1 >>
rect 128 38 129 39 
<< m1 >>
rect 13 39 14 40 
<< m1 >>
rect 19 39 20 40 
<< m2 >>
rect 19 39 20 40 
<< m1 >>
rect 51 39 52 40 
<< m2 >>
rect 51 39 52 40 
<< m2c >>
rect 51 39 52 40 
<< m1 >>
rect 51 39 52 40 
<< m2 >>
rect 51 39 52 40 
<< m2 >>
rect 52 39 53 40 
<< m1 >>
rect 53 39 54 40 
<< m2 >>
rect 53 39 54 40 
<< m1 >>
rect 54 39 55 40 
<< m2 >>
rect 54 39 55 40 
<< m1 >>
rect 55 39 56 40 
<< m2 >>
rect 55 39 56 40 
<< m1 >>
rect 56 39 57 40 
<< m1 >>
rect 57 39 58 40 
<< m1 >>
rect 58 39 59 40 
<< m1 >>
rect 59 39 60 40 
<< m1 >>
rect 60 39 61 40 
<< m1 >>
rect 61 39 62 40 
<< m1 >>
rect 62 39 63 40 
<< m1 >>
rect 63 39 64 40 
<< m1 >>
rect 64 39 65 40 
<< m1 >>
rect 68 39 69 40 
<< m2 >>
rect 68 39 69 40 
<< m2c >>
rect 68 39 69 40 
<< m1 >>
rect 68 39 69 40 
<< m2 >>
rect 68 39 69 40 
<< m1 >>
rect 69 39 70 40 
<< m1 >>
rect 70 39 71 40 
<< m1 >>
rect 71 39 72 40 
<< m1 >>
rect 72 39 73 40 
<< m1 >>
rect 73 39 74 40 
<< m1 >>
rect 86 39 87 40 
<< m2 >>
rect 86 39 87 40 
<< m2c >>
rect 86 39 87 40 
<< m1 >>
rect 86 39 87 40 
<< m2 >>
rect 86 39 87 40 
<< m1 >>
rect 87 39 88 40 
<< m1 >>
rect 88 39 89 40 
<< m1 >>
rect 89 39 90 40 
<< m2 >>
rect 89 39 90 40 
<< m2c >>
rect 89 39 90 40 
<< m1 >>
rect 89 39 90 40 
<< m2 >>
rect 89 39 90 40 
<< m2 >>
rect 90 39 91 40 
<< m1 >>
rect 91 39 92 40 
<< m2 >>
rect 91 39 92 40 
<< m2 >>
rect 92 39 93 40 
<< m1 >>
rect 93 39 94 40 
<< m2 >>
rect 93 39 94 40 
<< m2c >>
rect 93 39 94 40 
<< m1 >>
rect 93 39 94 40 
<< m2 >>
rect 93 39 94 40 
<< m1 >>
rect 94 39 95 40 
<< m1 >>
rect 95 39 96 40 
<< m2 >>
rect 95 39 96 40 
<< m2c >>
rect 95 39 96 40 
<< m1 >>
rect 95 39 96 40 
<< m2 >>
rect 95 39 96 40 
<< m1 >>
rect 100 39 101 40 
<< m1 >>
rect 121 39 122 40 
<< m1 >>
rect 128 39 129 40 
<< m2 >>
rect 128 39 129 40 
<< m2c >>
rect 128 39 129 40 
<< m1 >>
rect 128 39 129 40 
<< m2 >>
rect 128 39 129 40 
<< m1 >>
rect 13 40 14 41 
<< m1 >>
rect 19 40 20 41 
<< m2 >>
rect 19 40 20 41 
<< m1 >>
rect 20 40 21 41 
<< m2 >>
rect 20 40 21 41 
<< m1 >>
rect 21 40 22 41 
<< m2 >>
rect 21 40 22 41 
<< m1 >>
rect 22 40 23 41 
<< m2 >>
rect 22 40 23 41 
<< m1 >>
rect 23 40 24 41 
<< m2 >>
rect 23 40 24 41 
<< m1 >>
rect 24 40 25 41 
<< m2 >>
rect 24 40 25 41 
<< m1 >>
rect 25 40 26 41 
<< m2 >>
rect 25 40 26 41 
<< m1 >>
rect 26 40 27 41 
<< m2 >>
rect 26 40 27 41 
<< m1 >>
rect 27 40 28 41 
<< m2 >>
rect 27 40 28 41 
<< m1 >>
rect 28 40 29 41 
<< m2 >>
rect 28 40 29 41 
<< m1 >>
rect 29 40 30 41 
<< m2 >>
rect 29 40 30 41 
<< m1 >>
rect 30 40 31 41 
<< m2 >>
rect 30 40 31 41 
<< m1 >>
rect 31 40 32 41 
<< m2 >>
rect 31 40 32 41 
<< m1 >>
rect 32 40 33 41 
<< m2 >>
rect 32 40 33 41 
<< m1 >>
rect 33 40 34 41 
<< m2 >>
rect 33 40 34 41 
<< m1 >>
rect 34 40 35 41 
<< m2 >>
rect 34 40 35 41 
<< m1 >>
rect 35 40 36 41 
<< m2 >>
rect 35 40 36 41 
<< m1 >>
rect 36 40 37 41 
<< m2 >>
rect 36 40 37 41 
<< m1 >>
rect 37 40 38 41 
<< m2 >>
rect 37 40 38 41 
<< m2 >>
rect 38 40 39 41 
<< m1 >>
rect 39 40 40 41 
<< m2 >>
rect 39 40 40 41 
<< m2c >>
rect 39 40 40 41 
<< m1 >>
rect 39 40 40 41 
<< m2 >>
rect 39 40 40 41 
<< m1 >>
rect 51 40 52 41 
<< m1 >>
rect 53 40 54 41 
<< m2 >>
rect 68 40 69 41 
<< m2 >>
rect 86 40 87 41 
<< m1 >>
rect 91 40 92 41 
<< m2 >>
rect 95 40 96 41 
<< m1 >>
rect 100 40 101 41 
<< m1 >>
rect 121 40 122 41 
<< m2 >>
rect 128 40 129 41 
<< m1 >>
rect 13 41 14 42 
<< m1 >>
rect 37 41 38 42 
<< m1 >>
rect 39 41 40 42 
<< m1 >>
rect 51 41 52 42 
<< m1 >>
rect 53 41 54 42 
<< m1 >>
rect 55 41 56 42 
<< m1 >>
rect 56 41 57 42 
<< m1 >>
rect 57 41 58 42 
<< m1 >>
rect 58 41 59 42 
<< m1 >>
rect 59 41 60 42 
<< m1 >>
rect 60 41 61 42 
<< m1 >>
rect 61 41 62 42 
<< m1 >>
rect 62 41 63 42 
<< m1 >>
rect 63 41 64 42 
<< m1 >>
rect 64 41 65 42 
<< m1 >>
rect 65 41 66 42 
<< m1 >>
rect 66 41 67 42 
<< m1 >>
rect 67 41 68 42 
<< m1 >>
rect 68 41 69 42 
<< m2 >>
rect 68 41 69 42 
<< m1 >>
rect 69 41 70 42 
<< m1 >>
rect 70 41 71 42 
<< m1 >>
rect 71 41 72 42 
<< m1 >>
rect 72 41 73 42 
<< m1 >>
rect 73 41 74 42 
<< m1 >>
rect 74 41 75 42 
<< m1 >>
rect 75 41 76 42 
<< m1 >>
rect 76 41 77 42 
<< m1 >>
rect 77 41 78 42 
<< m1 >>
rect 78 41 79 42 
<< m1 >>
rect 79 41 80 42 
<< m1 >>
rect 80 41 81 42 
<< m1 >>
rect 81 41 82 42 
<< m1 >>
rect 82 41 83 42 
<< m1 >>
rect 83 41 84 42 
<< m1 >>
rect 84 41 85 42 
<< m1 >>
rect 85 41 86 42 
<< m1 >>
rect 86 41 87 42 
<< m2 >>
rect 86 41 87 42 
<< m1 >>
rect 87 41 88 42 
<< m1 >>
rect 88 41 89 42 
<< m1 >>
rect 89 41 90 42 
<< m2 >>
rect 89 41 90 42 
<< m2c >>
rect 89 41 90 42 
<< m1 >>
rect 89 41 90 42 
<< m2 >>
rect 89 41 90 42 
<< m2 >>
rect 90 41 91 42 
<< m1 >>
rect 91 41 92 42 
<< m2 >>
rect 91 41 92 42 
<< m2 >>
rect 92 41 93 42 
<< m1 >>
rect 93 41 94 42 
<< m2 >>
rect 93 41 94 42 
<< m2c >>
rect 93 41 94 42 
<< m1 >>
rect 93 41 94 42 
<< m2 >>
rect 93 41 94 42 
<< m1 >>
rect 94 41 95 42 
<< m1 >>
rect 95 41 96 42 
<< m2 >>
rect 95 41 96 42 
<< m1 >>
rect 96 41 97 42 
<< m1 >>
rect 97 41 98 42 
<< m1 >>
rect 98 41 99 42 
<< m2 >>
rect 98 41 99 42 
<< m2c >>
rect 98 41 99 42 
<< m1 >>
rect 98 41 99 42 
<< m2 >>
rect 98 41 99 42 
<< m2 >>
rect 99 41 100 42 
<< m1 >>
rect 100 41 101 42 
<< m2 >>
rect 100 41 101 42 
<< m2 >>
rect 101 41 102 42 
<< m1 >>
rect 102 41 103 42 
<< m2 >>
rect 102 41 103 42 
<< m2c >>
rect 102 41 103 42 
<< m1 >>
rect 102 41 103 42 
<< m2 >>
rect 102 41 103 42 
<< m1 >>
rect 103 41 104 42 
<< m1 >>
rect 104 41 105 42 
<< m1 >>
rect 105 41 106 42 
<< m1 >>
rect 106 41 107 42 
<< m1 >>
rect 107 41 108 42 
<< m1 >>
rect 108 41 109 42 
<< m1 >>
rect 109 41 110 42 
<< m1 >>
rect 110 41 111 42 
<< m1 >>
rect 111 41 112 42 
<< m1 >>
rect 112 41 113 42 
<< m1 >>
rect 113 41 114 42 
<< m1 >>
rect 114 41 115 42 
<< m1 >>
rect 115 41 116 42 
<< m1 >>
rect 116 41 117 42 
<< m1 >>
rect 117 41 118 42 
<< m1 >>
rect 118 41 119 42 
<< m1 >>
rect 119 41 120 42 
<< m2 >>
rect 119 41 120 42 
<< m2c >>
rect 119 41 120 42 
<< m1 >>
rect 119 41 120 42 
<< m2 >>
rect 119 41 120 42 
<< m2 >>
rect 120 41 121 42 
<< m1 >>
rect 121 41 122 42 
<< m2 >>
rect 121 41 122 42 
<< m2 >>
rect 122 41 123 42 
<< m1 >>
rect 123 41 124 42 
<< m2 >>
rect 123 41 124 42 
<< m2c >>
rect 123 41 124 42 
<< m1 >>
rect 123 41 124 42 
<< m2 >>
rect 123 41 124 42 
<< m1 >>
rect 124 41 125 42 
<< m1 >>
rect 125 41 126 42 
<< m1 >>
rect 126 41 127 42 
<< m1 >>
rect 127 41 128 42 
<< m1 >>
rect 128 41 129 42 
<< m2 >>
rect 128 41 129 42 
<< m1 >>
rect 129 41 130 42 
<< m1 >>
rect 130 41 131 42 
<< m1 >>
rect 131 41 132 42 
<< m1 >>
rect 132 41 133 42 
<< m1 >>
rect 133 41 134 42 
<< m1 >>
rect 134 41 135 42 
<< m1 >>
rect 135 41 136 42 
<< m1 >>
rect 13 42 14 43 
<< m1 >>
rect 14 42 15 43 
<< m1 >>
rect 15 42 16 43 
<< m1 >>
rect 16 42 17 43 
<< m1 >>
rect 17 42 18 43 
<< m1 >>
rect 18 42 19 43 
<< m1 >>
rect 19 42 20 43 
<< m1 >>
rect 20 42 21 43 
<< m1 >>
rect 21 42 22 43 
<< m1 >>
rect 22 42 23 43 
<< m1 >>
rect 23 42 24 43 
<< m1 >>
rect 24 42 25 43 
<< m1 >>
rect 25 42 26 43 
<< m1 >>
rect 26 42 27 43 
<< m1 >>
rect 27 42 28 43 
<< m1 >>
rect 28 42 29 43 
<< m1 >>
rect 29 42 30 43 
<< m1 >>
rect 30 42 31 43 
<< m1 >>
rect 31 42 32 43 
<< m1 >>
rect 32 42 33 43 
<< m1 >>
rect 33 42 34 43 
<< m1 >>
rect 34 42 35 43 
<< m1 >>
rect 35 42 36 43 
<< m2 >>
rect 35 42 36 43 
<< m2c >>
rect 35 42 36 43 
<< m1 >>
rect 35 42 36 43 
<< m2 >>
rect 35 42 36 43 
<< m2 >>
rect 36 42 37 43 
<< m1 >>
rect 37 42 38 43 
<< m2 >>
rect 37 42 38 43 
<< m2 >>
rect 38 42 39 43 
<< m1 >>
rect 39 42 40 43 
<< m2 >>
rect 39 42 40 43 
<< m2 >>
rect 40 42 41 43 
<< m1 >>
rect 41 42 42 43 
<< m2 >>
rect 41 42 42 43 
<< m2c >>
rect 41 42 42 43 
<< m1 >>
rect 41 42 42 43 
<< m2 >>
rect 41 42 42 43 
<< m1 >>
rect 42 42 43 43 
<< m1 >>
rect 43 42 44 43 
<< m1 >>
rect 44 42 45 43 
<< m1 >>
rect 45 42 46 43 
<< m1 >>
rect 46 42 47 43 
<< m1 >>
rect 47 42 48 43 
<< m1 >>
rect 48 42 49 43 
<< m1 >>
rect 49 42 50 43 
<< m1 >>
rect 50 42 51 43 
<< m1 >>
rect 51 42 52 43 
<< m1 >>
rect 53 42 54 43 
<< m1 >>
rect 55 42 56 43 
<< m2 >>
rect 68 42 69 43 
<< m2 >>
rect 70 42 71 43 
<< m2 >>
rect 71 42 72 43 
<< m2 >>
rect 72 42 73 43 
<< m2 >>
rect 73 42 74 43 
<< m2 >>
rect 74 42 75 43 
<< m2 >>
rect 75 42 76 43 
<< m2 >>
rect 76 42 77 43 
<< m2 >>
rect 77 42 78 43 
<< m2 >>
rect 78 42 79 43 
<< m2 >>
rect 79 42 80 43 
<< m2 >>
rect 80 42 81 43 
<< m2 >>
rect 81 42 82 43 
<< m2 >>
rect 82 42 83 43 
<< m2 >>
rect 83 42 84 43 
<< m2 >>
rect 84 42 85 43 
<< m2 >>
rect 85 42 86 43 
<< m2 >>
rect 86 42 87 43 
<< m1 >>
rect 91 42 92 43 
<< m2 >>
rect 95 42 96 43 
<< m1 >>
rect 100 42 101 43 
<< m1 >>
rect 121 42 122 43 
<< m2 >>
rect 128 42 129 43 
<< m1 >>
rect 135 42 136 43 
<< m1 >>
rect 37 43 38 44 
<< m1 >>
rect 39 43 40 44 
<< m1 >>
rect 53 43 54 44 
<< m2 >>
rect 53 43 54 44 
<< m2c >>
rect 53 43 54 44 
<< m1 >>
rect 53 43 54 44 
<< m2 >>
rect 53 43 54 44 
<< m1 >>
rect 55 43 56 44 
<< m2 >>
rect 55 43 56 44 
<< m2c >>
rect 55 43 56 44 
<< m1 >>
rect 55 43 56 44 
<< m2 >>
rect 55 43 56 44 
<< m1 >>
rect 68 43 69 44 
<< m2 >>
rect 68 43 69 44 
<< m2c >>
rect 68 43 69 44 
<< m1 >>
rect 68 43 69 44 
<< m2 >>
rect 68 43 69 44 
<< m1 >>
rect 70 43 71 44 
<< m2 >>
rect 70 43 71 44 
<< m2c >>
rect 70 43 71 44 
<< m1 >>
rect 70 43 71 44 
<< m2 >>
rect 70 43 71 44 
<< m1 >>
rect 91 43 92 44 
<< m2 >>
rect 91 43 92 44 
<< m2c >>
rect 91 43 92 44 
<< m1 >>
rect 91 43 92 44 
<< m2 >>
rect 91 43 92 44 
<< m1 >>
rect 95 43 96 44 
<< m2 >>
rect 95 43 96 44 
<< m2c >>
rect 95 43 96 44 
<< m1 >>
rect 95 43 96 44 
<< m2 >>
rect 95 43 96 44 
<< m1 >>
rect 96 43 97 44 
<< m1 >>
rect 97 43 98 44 
<< m1 >>
rect 98 43 99 44 
<< m2 >>
rect 98 43 99 44 
<< m2c >>
rect 98 43 99 44 
<< m1 >>
rect 98 43 99 44 
<< m2 >>
rect 98 43 99 44 
<< m2 >>
rect 99 43 100 44 
<< m1 >>
rect 100 43 101 44 
<< m2 >>
rect 100 43 101 44 
<< m2 >>
rect 101 43 102 44 
<< m1 >>
rect 102 43 103 44 
<< m2 >>
rect 102 43 103 44 
<< m2c >>
rect 102 43 103 44 
<< m1 >>
rect 102 43 103 44 
<< m2 >>
rect 102 43 103 44 
<< m1 >>
rect 103 43 104 44 
<< m1 >>
rect 109 43 110 44 
<< m2 >>
rect 109 43 110 44 
<< m1 >>
rect 110 43 111 44 
<< m2 >>
rect 110 43 111 44 
<< m1 >>
rect 111 43 112 44 
<< m2 >>
rect 111 43 112 44 
<< m1 >>
rect 112 43 113 44 
<< m2 >>
rect 112 43 113 44 
<< m1 >>
rect 113 43 114 44 
<< m2 >>
rect 113 43 114 44 
<< m1 >>
rect 114 43 115 44 
<< m2 >>
rect 114 43 115 44 
<< m1 >>
rect 115 43 116 44 
<< m2 >>
rect 115 43 116 44 
<< m1 >>
rect 116 43 117 44 
<< m2 >>
rect 116 43 117 44 
<< m1 >>
rect 117 43 118 44 
<< m2 >>
rect 117 43 118 44 
<< m1 >>
rect 118 43 119 44 
<< m2 >>
rect 118 43 119 44 
<< m1 >>
rect 119 43 120 44 
<< m2 >>
rect 119 43 120 44 
<< m1 >>
rect 120 43 121 44 
<< m2 >>
rect 120 43 121 44 
<< m1 >>
rect 121 43 122 44 
<< m2 >>
rect 121 43 122 44 
<< m2 >>
rect 122 43 123 44 
<< m1 >>
rect 123 43 124 44 
<< m2 >>
rect 123 43 124 44 
<< m2c >>
rect 123 43 124 44 
<< m1 >>
rect 123 43 124 44 
<< m2 >>
rect 123 43 124 44 
<< m1 >>
rect 124 43 125 44 
<< m1 >>
rect 128 43 129 44 
<< m2 >>
rect 128 43 129 44 
<< m2c >>
rect 128 43 129 44 
<< m1 >>
rect 128 43 129 44 
<< m2 >>
rect 128 43 129 44 
<< m1 >>
rect 135 43 136 44 
<< m1 >>
rect 37 44 38 45 
<< m1 >>
rect 39 44 40 45 
<< m2 >>
rect 52 44 53 45 
<< m2 >>
rect 53 44 54 45 
<< m2 >>
rect 55 44 56 45 
<< m1 >>
rect 68 44 69 45 
<< m1 >>
rect 70 44 71 45 
<< m2 >>
rect 91 44 92 45 
<< m1 >>
rect 100 44 101 45 
<< m1 >>
rect 103 44 104 45 
<< m1 >>
rect 109 44 110 45 
<< m2 >>
rect 109 44 110 45 
<< m1 >>
rect 124 44 125 45 
<< m1 >>
rect 128 44 129 45 
<< m1 >>
rect 135 44 136 45 
<< m2 >>
rect 135 44 136 45 
<< m2c >>
rect 135 44 136 45 
<< m1 >>
rect 135 44 136 45 
<< m2 >>
rect 135 44 136 45 
<< m1 >>
rect 37 45 38 46 
<< m1 >>
rect 39 45 40 46 
<< m1 >>
rect 49 45 50 46 
<< m1 >>
rect 50 45 51 46 
<< m1 >>
rect 51 45 52 46 
<< m1 >>
rect 52 45 53 46 
<< m2 >>
rect 52 45 53 46 
<< m1 >>
rect 53 45 54 46 
<< m1 >>
rect 54 45 55 46 
<< m1 >>
rect 55 45 56 46 
<< m2 >>
rect 55 45 56 46 
<< m1 >>
rect 56 45 57 46 
<< m1 >>
rect 57 45 58 46 
<< m1 >>
rect 58 45 59 46 
<< m1 >>
rect 59 45 60 46 
<< m1 >>
rect 60 45 61 46 
<< m1 >>
rect 61 45 62 46 
<< m1 >>
rect 62 45 63 46 
<< m1 >>
rect 63 45 64 46 
<< m1 >>
rect 64 45 65 46 
<< m1 >>
rect 68 45 69 46 
<< m2 >>
rect 68 45 69 46 
<< m2c >>
rect 68 45 69 46 
<< m1 >>
rect 68 45 69 46 
<< m2 >>
rect 68 45 69 46 
<< m2 >>
rect 69 45 70 46 
<< m1 >>
rect 70 45 71 46 
<< m2 >>
rect 70 45 71 46 
<< m2 >>
rect 71 45 72 46 
<< m1 >>
rect 85 45 86 46 
<< m1 >>
rect 86 45 87 46 
<< m1 >>
rect 87 45 88 46 
<< m1 >>
rect 88 45 89 46 
<< m1 >>
rect 89 45 90 46 
<< m1 >>
rect 90 45 91 46 
<< m1 >>
rect 91 45 92 46 
<< m2 >>
rect 91 45 92 46 
<< m1 >>
rect 92 45 93 46 
<< m1 >>
rect 93 45 94 46 
<< m1 >>
rect 94 45 95 46 
<< m1 >>
rect 95 45 96 46 
<< m1 >>
rect 96 45 97 46 
<< m1 >>
rect 97 45 98 46 
<< m1 >>
rect 98 45 99 46 
<< m1 >>
rect 100 45 101 46 
<< m1 >>
rect 103 45 104 46 
<< m1 >>
rect 109 45 110 46 
<< m2 >>
rect 109 45 110 46 
<< m1 >>
rect 124 45 125 46 
<< m1 >>
rect 128 45 129 46 
<< m2 >>
rect 135 45 136 46 
<< m1 >>
rect 16 46 17 47 
<< m1 >>
rect 17 46 18 47 
<< m1 >>
rect 18 46 19 47 
<< m1 >>
rect 19 46 20 47 
<< m1 >>
rect 20 46 21 47 
<< m1 >>
rect 21 46 22 47 
<< m1 >>
rect 22 46 23 47 
<< m1 >>
rect 23 46 24 47 
<< m1 >>
rect 24 46 25 47 
<< m1 >>
rect 25 46 26 47 
<< m1 >>
rect 26 46 27 47 
<< m1 >>
rect 27 46 28 47 
<< m1 >>
rect 28 46 29 47 
<< m1 >>
rect 37 46 38 47 
<< m1 >>
rect 39 46 40 47 
<< m1 >>
rect 49 46 50 47 
<< m2 >>
rect 52 46 53 47 
<< m2 >>
rect 55 46 56 47 
<< m1 >>
rect 64 46 65 47 
<< m1 >>
rect 70 46 71 47 
<< m2 >>
rect 71 46 72 47 
<< m1 >>
rect 72 46 73 47 
<< m2 >>
rect 72 46 73 47 
<< m2c >>
rect 72 46 73 47 
<< m1 >>
rect 72 46 73 47 
<< m2 >>
rect 72 46 73 47 
<< m1 >>
rect 73 46 74 47 
<< m1 >>
rect 85 46 86 47 
<< m2 >>
rect 91 46 92 47 
<< m1 >>
rect 98 46 99 47 
<< m1 >>
rect 100 46 101 47 
<< m1 >>
rect 103 46 104 47 
<< m1 >>
rect 109 46 110 47 
<< m2 >>
rect 109 46 110 47 
<< m1 >>
rect 124 46 125 47 
<< m1 >>
rect 128 46 129 47 
<< m2 >>
rect 135 46 136 47 
<< m1 >>
rect 136 46 137 47 
<< m1 >>
rect 137 46 138 47 
<< m1 >>
rect 138 46 139 47 
<< m1 >>
rect 139 46 140 47 
<< m1 >>
rect 142 46 143 47 
<< m1 >>
rect 143 46 144 47 
<< m1 >>
rect 144 46 145 47 
<< m1 >>
rect 145 46 146 47 
<< m1 >>
rect 16 47 17 48 
<< m1 >>
rect 28 47 29 48 
<< m1 >>
rect 37 47 38 48 
<< m1 >>
rect 39 47 40 48 
<< m1 >>
rect 49 47 50 48 
<< m1 >>
rect 52 47 53 48 
<< m2 >>
rect 52 47 53 48 
<< m2c >>
rect 52 47 53 48 
<< m1 >>
rect 52 47 53 48 
<< m2 >>
rect 52 47 53 48 
<< m1 >>
rect 55 47 56 48 
<< m2 >>
rect 55 47 56 48 
<< m2c >>
rect 55 47 56 48 
<< m1 >>
rect 55 47 56 48 
<< m2 >>
rect 55 47 56 48 
<< m1 >>
rect 64 47 65 48 
<< m1 >>
rect 70 47 71 48 
<< m1 >>
rect 73 47 74 48 
<< m1 >>
rect 85 47 86 48 
<< m1 >>
rect 91 47 92 48 
<< m2 >>
rect 91 47 92 48 
<< m2c >>
rect 91 47 92 48 
<< m1 >>
rect 91 47 92 48 
<< m2 >>
rect 91 47 92 48 
<< m1 >>
rect 98 47 99 48 
<< m1 >>
rect 100 47 101 48 
<< m1 >>
rect 103 47 104 48 
<< m1 >>
rect 109 47 110 48 
<< m2 >>
rect 109 47 110 48 
<< m1 >>
rect 124 47 125 48 
<< m1 >>
rect 128 47 129 48 
<< m2 >>
rect 135 47 136 48 
<< m1 >>
rect 136 47 137 48 
<< m1 >>
rect 139 47 140 48 
<< m1 >>
rect 142 47 143 48 
<< m1 >>
rect 145 47 146 48 
<< pdiffusion >>
rect 12 48 13 49 
<< pdiffusion >>
rect 13 48 14 49 
<< pdiffusion >>
rect 14 48 15 49 
<< pdiffusion >>
rect 15 48 16 49 
<< m1 >>
rect 16 48 17 49 
<< pdiffusion >>
rect 16 48 17 49 
<< pdiffusion >>
rect 17 48 18 49 
<< m1 >>
rect 28 48 29 49 
<< pdiffusion >>
rect 30 48 31 49 
<< pdiffusion >>
rect 31 48 32 49 
<< pdiffusion >>
rect 32 48 33 49 
<< pdiffusion >>
rect 33 48 34 49 
<< pdiffusion >>
rect 34 48 35 49 
<< pdiffusion >>
rect 35 48 36 49 
<< m1 >>
rect 37 48 38 49 
<< m1 >>
rect 39 48 40 49 
<< pdiffusion >>
rect 48 48 49 49 
<< m1 >>
rect 49 48 50 49 
<< pdiffusion >>
rect 49 48 50 49 
<< pdiffusion >>
rect 50 48 51 49 
<< pdiffusion >>
rect 51 48 52 49 
<< m1 >>
rect 52 48 53 49 
<< pdiffusion >>
rect 52 48 53 49 
<< pdiffusion >>
rect 53 48 54 49 
<< m1 >>
rect 55 48 56 49 
<< m1 >>
rect 64 48 65 49 
<< pdiffusion >>
rect 66 48 67 49 
<< pdiffusion >>
rect 67 48 68 49 
<< pdiffusion >>
rect 68 48 69 49 
<< pdiffusion >>
rect 69 48 70 49 
<< m1 >>
rect 70 48 71 49 
<< pdiffusion >>
rect 70 48 71 49 
<< pdiffusion >>
rect 71 48 72 49 
<< m1 >>
rect 73 48 74 49 
<< pdiffusion >>
rect 84 48 85 49 
<< m1 >>
rect 85 48 86 49 
<< pdiffusion >>
rect 85 48 86 49 
<< pdiffusion >>
rect 86 48 87 49 
<< pdiffusion >>
rect 87 48 88 49 
<< pdiffusion >>
rect 88 48 89 49 
<< pdiffusion >>
rect 89 48 90 49 
<< m1 >>
rect 91 48 92 49 
<< m1 >>
rect 98 48 99 49 
<< m1 >>
rect 100 48 101 49 
<< pdiffusion >>
rect 102 48 103 49 
<< m1 >>
rect 103 48 104 49 
<< pdiffusion >>
rect 103 48 104 49 
<< pdiffusion >>
rect 104 48 105 49 
<< pdiffusion >>
rect 105 48 106 49 
<< pdiffusion >>
rect 106 48 107 49 
<< pdiffusion >>
rect 107 48 108 49 
<< m1 >>
rect 109 48 110 49 
<< m2 >>
rect 109 48 110 49 
<< pdiffusion >>
rect 120 48 121 49 
<< pdiffusion >>
rect 121 48 122 49 
<< pdiffusion >>
rect 122 48 123 49 
<< pdiffusion >>
rect 123 48 124 49 
<< m1 >>
rect 124 48 125 49 
<< pdiffusion >>
rect 124 48 125 49 
<< pdiffusion >>
rect 125 48 126 49 
<< m1 >>
rect 128 48 129 49 
<< m2 >>
rect 135 48 136 49 
<< m1 >>
rect 136 48 137 49 
<< pdiffusion >>
rect 138 48 139 49 
<< m1 >>
rect 139 48 140 49 
<< pdiffusion >>
rect 139 48 140 49 
<< pdiffusion >>
rect 140 48 141 49 
<< pdiffusion >>
rect 141 48 142 49 
<< m1 >>
rect 142 48 143 49 
<< pdiffusion >>
rect 142 48 143 49 
<< pdiffusion >>
rect 143 48 144 49 
<< m1 >>
rect 145 48 146 49 
<< pdiffusion >>
rect 12 49 13 50 
<< pdiffusion >>
rect 13 49 14 50 
<< pdiffusion >>
rect 14 49 15 50 
<< pdiffusion >>
rect 15 49 16 50 
<< pdiffusion >>
rect 16 49 17 50 
<< pdiffusion >>
rect 17 49 18 50 
<< m1 >>
rect 28 49 29 50 
<< pdiffusion >>
rect 30 49 31 50 
<< pdiffusion >>
rect 31 49 32 50 
<< pdiffusion >>
rect 32 49 33 50 
<< pdiffusion >>
rect 33 49 34 50 
<< pdiffusion >>
rect 34 49 35 50 
<< pdiffusion >>
rect 35 49 36 50 
<< m1 >>
rect 37 49 38 50 
<< m1 >>
rect 39 49 40 50 
<< pdiffusion >>
rect 48 49 49 50 
<< pdiffusion >>
rect 49 49 50 50 
<< pdiffusion >>
rect 50 49 51 50 
<< pdiffusion >>
rect 51 49 52 50 
<< pdiffusion >>
rect 52 49 53 50 
<< pdiffusion >>
rect 53 49 54 50 
<< m1 >>
rect 55 49 56 50 
<< m1 >>
rect 64 49 65 50 
<< pdiffusion >>
rect 66 49 67 50 
<< pdiffusion >>
rect 67 49 68 50 
<< pdiffusion >>
rect 68 49 69 50 
<< pdiffusion >>
rect 69 49 70 50 
<< pdiffusion >>
rect 70 49 71 50 
<< pdiffusion >>
rect 71 49 72 50 
<< m1 >>
rect 73 49 74 50 
<< pdiffusion >>
rect 84 49 85 50 
<< pdiffusion >>
rect 85 49 86 50 
<< pdiffusion >>
rect 86 49 87 50 
<< pdiffusion >>
rect 87 49 88 50 
<< pdiffusion >>
rect 88 49 89 50 
<< pdiffusion >>
rect 89 49 90 50 
<< m1 >>
rect 91 49 92 50 
<< m1 >>
rect 98 49 99 50 
<< m1 >>
rect 100 49 101 50 
<< pdiffusion >>
rect 102 49 103 50 
<< pdiffusion >>
rect 103 49 104 50 
<< pdiffusion >>
rect 104 49 105 50 
<< pdiffusion >>
rect 105 49 106 50 
<< pdiffusion >>
rect 106 49 107 50 
<< pdiffusion >>
rect 107 49 108 50 
<< m1 >>
rect 109 49 110 50 
<< m2 >>
rect 109 49 110 50 
<< pdiffusion >>
rect 120 49 121 50 
<< pdiffusion >>
rect 121 49 122 50 
<< pdiffusion >>
rect 122 49 123 50 
<< pdiffusion >>
rect 123 49 124 50 
<< pdiffusion >>
rect 124 49 125 50 
<< pdiffusion >>
rect 125 49 126 50 
<< m1 >>
rect 128 49 129 50 
<< m2 >>
rect 135 49 136 50 
<< m1 >>
rect 136 49 137 50 
<< pdiffusion >>
rect 138 49 139 50 
<< pdiffusion >>
rect 139 49 140 50 
<< pdiffusion >>
rect 140 49 141 50 
<< pdiffusion >>
rect 141 49 142 50 
<< pdiffusion >>
rect 142 49 143 50 
<< pdiffusion >>
rect 143 49 144 50 
<< m1 >>
rect 145 49 146 50 
<< pdiffusion >>
rect 12 50 13 51 
<< pdiffusion >>
rect 13 50 14 51 
<< pdiffusion >>
rect 14 50 15 51 
<< pdiffusion >>
rect 15 50 16 51 
<< pdiffusion >>
rect 16 50 17 51 
<< pdiffusion >>
rect 17 50 18 51 
<< m1 >>
rect 28 50 29 51 
<< pdiffusion >>
rect 30 50 31 51 
<< pdiffusion >>
rect 31 50 32 51 
<< pdiffusion >>
rect 32 50 33 51 
<< pdiffusion >>
rect 33 50 34 51 
<< pdiffusion >>
rect 34 50 35 51 
<< pdiffusion >>
rect 35 50 36 51 
<< m1 >>
rect 37 50 38 51 
<< m1 >>
rect 39 50 40 51 
<< pdiffusion >>
rect 48 50 49 51 
<< pdiffusion >>
rect 49 50 50 51 
<< pdiffusion >>
rect 50 50 51 51 
<< pdiffusion >>
rect 51 50 52 51 
<< pdiffusion >>
rect 52 50 53 51 
<< pdiffusion >>
rect 53 50 54 51 
<< m1 >>
rect 55 50 56 51 
<< m1 >>
rect 64 50 65 51 
<< pdiffusion >>
rect 66 50 67 51 
<< pdiffusion >>
rect 67 50 68 51 
<< pdiffusion >>
rect 68 50 69 51 
<< pdiffusion >>
rect 69 50 70 51 
<< pdiffusion >>
rect 70 50 71 51 
<< pdiffusion >>
rect 71 50 72 51 
<< m1 >>
rect 73 50 74 51 
<< pdiffusion >>
rect 84 50 85 51 
<< pdiffusion >>
rect 85 50 86 51 
<< pdiffusion >>
rect 86 50 87 51 
<< pdiffusion >>
rect 87 50 88 51 
<< pdiffusion >>
rect 88 50 89 51 
<< pdiffusion >>
rect 89 50 90 51 
<< m1 >>
rect 91 50 92 51 
<< m1 >>
rect 98 50 99 51 
<< m1 >>
rect 100 50 101 51 
<< pdiffusion >>
rect 102 50 103 51 
<< pdiffusion >>
rect 103 50 104 51 
<< pdiffusion >>
rect 104 50 105 51 
<< pdiffusion >>
rect 105 50 106 51 
<< pdiffusion >>
rect 106 50 107 51 
<< pdiffusion >>
rect 107 50 108 51 
<< m1 >>
rect 109 50 110 51 
<< m2 >>
rect 109 50 110 51 
<< pdiffusion >>
rect 120 50 121 51 
<< pdiffusion >>
rect 121 50 122 51 
<< pdiffusion >>
rect 122 50 123 51 
<< pdiffusion >>
rect 123 50 124 51 
<< pdiffusion >>
rect 124 50 125 51 
<< pdiffusion >>
rect 125 50 126 51 
<< m1 >>
rect 128 50 129 51 
<< m2 >>
rect 135 50 136 51 
<< m1 >>
rect 136 50 137 51 
<< pdiffusion >>
rect 138 50 139 51 
<< pdiffusion >>
rect 139 50 140 51 
<< pdiffusion >>
rect 140 50 141 51 
<< pdiffusion >>
rect 141 50 142 51 
<< pdiffusion >>
rect 142 50 143 51 
<< pdiffusion >>
rect 143 50 144 51 
<< m1 >>
rect 145 50 146 51 
<< pdiffusion >>
rect 12 51 13 52 
<< pdiffusion >>
rect 13 51 14 52 
<< pdiffusion >>
rect 14 51 15 52 
<< pdiffusion >>
rect 15 51 16 52 
<< pdiffusion >>
rect 16 51 17 52 
<< pdiffusion >>
rect 17 51 18 52 
<< m1 >>
rect 28 51 29 52 
<< pdiffusion >>
rect 30 51 31 52 
<< pdiffusion >>
rect 31 51 32 52 
<< pdiffusion >>
rect 32 51 33 52 
<< pdiffusion >>
rect 33 51 34 52 
<< pdiffusion >>
rect 34 51 35 52 
<< pdiffusion >>
rect 35 51 36 52 
<< m1 >>
rect 37 51 38 52 
<< m1 >>
rect 39 51 40 52 
<< pdiffusion >>
rect 48 51 49 52 
<< pdiffusion >>
rect 49 51 50 52 
<< pdiffusion >>
rect 50 51 51 52 
<< pdiffusion >>
rect 51 51 52 52 
<< pdiffusion >>
rect 52 51 53 52 
<< pdiffusion >>
rect 53 51 54 52 
<< m1 >>
rect 55 51 56 52 
<< m1 >>
rect 64 51 65 52 
<< pdiffusion >>
rect 66 51 67 52 
<< pdiffusion >>
rect 67 51 68 52 
<< pdiffusion >>
rect 68 51 69 52 
<< pdiffusion >>
rect 69 51 70 52 
<< pdiffusion >>
rect 70 51 71 52 
<< pdiffusion >>
rect 71 51 72 52 
<< m1 >>
rect 73 51 74 52 
<< pdiffusion >>
rect 84 51 85 52 
<< pdiffusion >>
rect 85 51 86 52 
<< pdiffusion >>
rect 86 51 87 52 
<< pdiffusion >>
rect 87 51 88 52 
<< pdiffusion >>
rect 88 51 89 52 
<< pdiffusion >>
rect 89 51 90 52 
<< m1 >>
rect 91 51 92 52 
<< m1 >>
rect 98 51 99 52 
<< m1 >>
rect 100 51 101 52 
<< pdiffusion >>
rect 102 51 103 52 
<< pdiffusion >>
rect 103 51 104 52 
<< pdiffusion >>
rect 104 51 105 52 
<< pdiffusion >>
rect 105 51 106 52 
<< pdiffusion >>
rect 106 51 107 52 
<< pdiffusion >>
rect 107 51 108 52 
<< m1 >>
rect 109 51 110 52 
<< m2 >>
rect 109 51 110 52 
<< pdiffusion >>
rect 120 51 121 52 
<< pdiffusion >>
rect 121 51 122 52 
<< pdiffusion >>
rect 122 51 123 52 
<< pdiffusion >>
rect 123 51 124 52 
<< pdiffusion >>
rect 124 51 125 52 
<< pdiffusion >>
rect 125 51 126 52 
<< m1 >>
rect 128 51 129 52 
<< m2 >>
rect 135 51 136 52 
<< m1 >>
rect 136 51 137 52 
<< pdiffusion >>
rect 138 51 139 52 
<< pdiffusion >>
rect 139 51 140 52 
<< pdiffusion >>
rect 140 51 141 52 
<< pdiffusion >>
rect 141 51 142 52 
<< pdiffusion >>
rect 142 51 143 52 
<< pdiffusion >>
rect 143 51 144 52 
<< m1 >>
rect 145 51 146 52 
<< pdiffusion >>
rect 12 52 13 53 
<< pdiffusion >>
rect 13 52 14 53 
<< pdiffusion >>
rect 14 52 15 53 
<< pdiffusion >>
rect 15 52 16 53 
<< pdiffusion >>
rect 16 52 17 53 
<< pdiffusion >>
rect 17 52 18 53 
<< m1 >>
rect 28 52 29 53 
<< pdiffusion >>
rect 30 52 31 53 
<< pdiffusion >>
rect 31 52 32 53 
<< pdiffusion >>
rect 32 52 33 53 
<< pdiffusion >>
rect 33 52 34 53 
<< pdiffusion >>
rect 34 52 35 53 
<< pdiffusion >>
rect 35 52 36 53 
<< m1 >>
rect 37 52 38 53 
<< m1 >>
rect 39 52 40 53 
<< pdiffusion >>
rect 48 52 49 53 
<< pdiffusion >>
rect 49 52 50 53 
<< pdiffusion >>
rect 50 52 51 53 
<< pdiffusion >>
rect 51 52 52 53 
<< pdiffusion >>
rect 52 52 53 53 
<< pdiffusion >>
rect 53 52 54 53 
<< m1 >>
rect 55 52 56 53 
<< m1 >>
rect 64 52 65 53 
<< pdiffusion >>
rect 66 52 67 53 
<< pdiffusion >>
rect 67 52 68 53 
<< pdiffusion >>
rect 68 52 69 53 
<< pdiffusion >>
rect 69 52 70 53 
<< pdiffusion >>
rect 70 52 71 53 
<< pdiffusion >>
rect 71 52 72 53 
<< m1 >>
rect 73 52 74 53 
<< pdiffusion >>
rect 84 52 85 53 
<< pdiffusion >>
rect 85 52 86 53 
<< pdiffusion >>
rect 86 52 87 53 
<< pdiffusion >>
rect 87 52 88 53 
<< pdiffusion >>
rect 88 52 89 53 
<< pdiffusion >>
rect 89 52 90 53 
<< m1 >>
rect 91 52 92 53 
<< m1 >>
rect 98 52 99 53 
<< m1 >>
rect 100 52 101 53 
<< pdiffusion >>
rect 102 52 103 53 
<< pdiffusion >>
rect 103 52 104 53 
<< pdiffusion >>
rect 104 52 105 53 
<< pdiffusion >>
rect 105 52 106 53 
<< pdiffusion >>
rect 106 52 107 53 
<< pdiffusion >>
rect 107 52 108 53 
<< m1 >>
rect 109 52 110 53 
<< m2 >>
rect 109 52 110 53 
<< pdiffusion >>
rect 120 52 121 53 
<< pdiffusion >>
rect 121 52 122 53 
<< pdiffusion >>
rect 122 52 123 53 
<< pdiffusion >>
rect 123 52 124 53 
<< pdiffusion >>
rect 124 52 125 53 
<< pdiffusion >>
rect 125 52 126 53 
<< m1 >>
rect 128 52 129 53 
<< m2 >>
rect 135 52 136 53 
<< m1 >>
rect 136 52 137 53 
<< pdiffusion >>
rect 138 52 139 53 
<< pdiffusion >>
rect 139 52 140 53 
<< pdiffusion >>
rect 140 52 141 53 
<< pdiffusion >>
rect 141 52 142 53 
<< pdiffusion >>
rect 142 52 143 53 
<< pdiffusion >>
rect 143 52 144 53 
<< m1 >>
rect 145 52 146 53 
<< pdiffusion >>
rect 12 53 13 54 
<< m1 >>
rect 13 53 14 54 
<< pdiffusion >>
rect 13 53 14 54 
<< pdiffusion >>
rect 14 53 15 54 
<< pdiffusion >>
rect 15 53 16 54 
<< m1 >>
rect 16 53 17 54 
<< pdiffusion >>
rect 16 53 17 54 
<< pdiffusion >>
rect 17 53 18 54 
<< m1 >>
rect 28 53 29 54 
<< pdiffusion >>
rect 30 53 31 54 
<< pdiffusion >>
rect 31 53 32 54 
<< pdiffusion >>
rect 32 53 33 54 
<< pdiffusion >>
rect 33 53 34 54 
<< m1 >>
rect 34 53 35 54 
<< pdiffusion >>
rect 34 53 35 54 
<< pdiffusion >>
rect 35 53 36 54 
<< m1 >>
rect 37 53 38 54 
<< m1 >>
rect 39 53 40 54 
<< pdiffusion >>
rect 48 53 49 54 
<< m1 >>
rect 49 53 50 54 
<< pdiffusion >>
rect 49 53 50 54 
<< pdiffusion >>
rect 50 53 51 54 
<< pdiffusion >>
rect 51 53 52 54 
<< m1 >>
rect 52 53 53 54 
<< pdiffusion >>
rect 52 53 53 54 
<< pdiffusion >>
rect 53 53 54 54 
<< m1 >>
rect 55 53 56 54 
<< m1 >>
rect 64 53 65 54 
<< pdiffusion >>
rect 66 53 67 54 
<< m1 >>
rect 67 53 68 54 
<< pdiffusion >>
rect 67 53 68 54 
<< pdiffusion >>
rect 68 53 69 54 
<< pdiffusion >>
rect 69 53 70 54 
<< pdiffusion >>
rect 70 53 71 54 
<< pdiffusion >>
rect 71 53 72 54 
<< m1 >>
rect 73 53 74 54 
<< pdiffusion >>
rect 84 53 85 54 
<< m1 >>
rect 85 53 86 54 
<< pdiffusion >>
rect 85 53 86 54 
<< pdiffusion >>
rect 86 53 87 54 
<< pdiffusion >>
rect 87 53 88 54 
<< pdiffusion >>
rect 88 53 89 54 
<< pdiffusion >>
rect 89 53 90 54 
<< m1 >>
rect 91 53 92 54 
<< m1 >>
rect 98 53 99 54 
<< m1 >>
rect 100 53 101 54 
<< pdiffusion >>
rect 102 53 103 54 
<< pdiffusion >>
rect 103 53 104 54 
<< pdiffusion >>
rect 104 53 105 54 
<< pdiffusion >>
rect 105 53 106 54 
<< m1 >>
rect 106 53 107 54 
<< pdiffusion >>
rect 106 53 107 54 
<< pdiffusion >>
rect 107 53 108 54 
<< m1 >>
rect 109 53 110 54 
<< m2 >>
rect 109 53 110 54 
<< pdiffusion >>
rect 120 53 121 54 
<< m1 >>
rect 121 53 122 54 
<< pdiffusion >>
rect 121 53 122 54 
<< pdiffusion >>
rect 122 53 123 54 
<< pdiffusion >>
rect 123 53 124 54 
<< pdiffusion >>
rect 124 53 125 54 
<< pdiffusion >>
rect 125 53 126 54 
<< m1 >>
rect 128 53 129 54 
<< m2 >>
rect 135 53 136 54 
<< m1 >>
rect 136 53 137 54 
<< pdiffusion >>
rect 138 53 139 54 
<< pdiffusion >>
rect 139 53 140 54 
<< pdiffusion >>
rect 140 53 141 54 
<< pdiffusion >>
rect 141 53 142 54 
<< m1 >>
rect 142 53 143 54 
<< pdiffusion >>
rect 142 53 143 54 
<< pdiffusion >>
rect 143 53 144 54 
<< m1 >>
rect 145 53 146 54 
<< m1 >>
rect 13 54 14 55 
<< m1 >>
rect 16 54 17 55 
<< m1 >>
rect 28 54 29 55 
<< m1 >>
rect 34 54 35 55 
<< m1 >>
rect 37 54 38 55 
<< m1 >>
rect 39 54 40 55 
<< m1 >>
rect 49 54 50 55 
<< m1 >>
rect 52 54 53 55 
<< m1 >>
rect 55 54 56 55 
<< m1 >>
rect 64 54 65 55 
<< m1 >>
rect 67 54 68 55 
<< m1 >>
rect 73 54 74 55 
<< m1 >>
rect 85 54 86 55 
<< m1 >>
rect 91 54 92 55 
<< m1 >>
rect 98 54 99 55 
<< m1 >>
rect 100 54 101 55 
<< m1 >>
rect 106 54 107 55 
<< m1 >>
rect 109 54 110 55 
<< m2 >>
rect 109 54 110 55 
<< m1 >>
rect 121 54 122 55 
<< m1 >>
rect 128 54 129 55 
<< m2 >>
rect 135 54 136 55 
<< m1 >>
rect 136 54 137 55 
<< m1 >>
rect 142 54 143 55 
<< m1 >>
rect 145 54 146 55 
<< m1 >>
rect 13 55 14 56 
<< m1 >>
rect 16 55 17 56 
<< m1 >>
rect 28 55 29 56 
<< m1 >>
rect 34 55 35 56 
<< m1 >>
rect 37 55 38 56 
<< m1 >>
rect 39 55 40 56 
<< m1 >>
rect 40 55 41 56 
<< m1 >>
rect 41 55 42 56 
<< m1 >>
rect 42 55 43 56 
<< m1 >>
rect 43 55 44 56 
<< m1 >>
rect 44 55 45 56 
<< m1 >>
rect 45 55 46 56 
<< m1 >>
rect 46 55 47 56 
<< m1 >>
rect 47 55 48 56 
<< m1 >>
rect 48 55 49 56 
<< m1 >>
rect 49 55 50 56 
<< m1 >>
rect 52 55 53 56 
<< m1 >>
rect 55 55 56 56 
<< m1 >>
rect 64 55 65 56 
<< m1 >>
rect 67 55 68 56 
<< m1 >>
rect 73 55 74 56 
<< m1 >>
rect 85 55 86 56 
<< m1 >>
rect 91 55 92 56 
<< m1 >>
rect 98 55 99 56 
<< m1 >>
rect 100 55 101 56 
<< m1 >>
rect 106 55 107 56 
<< m1 >>
rect 107 55 108 56 
<< m1 >>
rect 108 55 109 56 
<< m1 >>
rect 109 55 110 56 
<< m2 >>
rect 109 55 110 56 
<< m1 >>
rect 121 55 122 56 
<< m1 >>
rect 128 55 129 56 
<< m2 >>
rect 135 55 136 56 
<< m1 >>
rect 136 55 137 56 
<< m2 >>
rect 136 55 137 56 
<< m2 >>
rect 137 55 138 56 
<< m1 >>
rect 138 55 139 56 
<< m2 >>
rect 138 55 139 56 
<< m2c >>
rect 138 55 139 56 
<< m1 >>
rect 138 55 139 56 
<< m2 >>
rect 138 55 139 56 
<< m1 >>
rect 142 55 143 56 
<< m1 >>
rect 145 55 146 56 
<< m1 >>
rect 13 56 14 57 
<< m1 >>
rect 16 56 17 57 
<< m1 >>
rect 28 56 29 57 
<< m1 >>
rect 29 56 30 57 
<< m1 >>
rect 30 56 31 57 
<< m2 >>
rect 30 56 31 57 
<< m2c >>
rect 30 56 31 57 
<< m1 >>
rect 30 56 31 57 
<< m2 >>
rect 30 56 31 57 
<< m1 >>
rect 34 56 35 57 
<< m2 >>
rect 34 56 35 57 
<< m2c >>
rect 34 56 35 57 
<< m1 >>
rect 34 56 35 57 
<< m2 >>
rect 34 56 35 57 
<< m1 >>
rect 37 56 38 57 
<< m2 >>
rect 37 56 38 57 
<< m2c >>
rect 37 56 38 57 
<< m1 >>
rect 37 56 38 57 
<< m2 >>
rect 37 56 38 57 
<< m1 >>
rect 52 56 53 57 
<< m2 >>
rect 52 56 53 57 
<< m2c >>
rect 52 56 53 57 
<< m1 >>
rect 52 56 53 57 
<< m2 >>
rect 52 56 53 57 
<< m1 >>
rect 55 56 56 57 
<< m2 >>
rect 55 56 56 57 
<< m2c >>
rect 55 56 56 57 
<< m1 >>
rect 55 56 56 57 
<< m2 >>
rect 55 56 56 57 
<< m1 >>
rect 57 56 58 57 
<< m2 >>
rect 57 56 58 57 
<< m2c >>
rect 57 56 58 57 
<< m1 >>
rect 57 56 58 57 
<< m2 >>
rect 57 56 58 57 
<< m1 >>
rect 58 56 59 57 
<< m1 >>
rect 59 56 60 57 
<< m1 >>
rect 60 56 61 57 
<< m1 >>
rect 61 56 62 57 
<< m1 >>
rect 62 56 63 57 
<< m2 >>
rect 62 56 63 57 
<< m2c >>
rect 62 56 63 57 
<< m1 >>
rect 62 56 63 57 
<< m2 >>
rect 62 56 63 57 
<< m2 >>
rect 63 56 64 57 
<< m1 >>
rect 64 56 65 57 
<< m2 >>
rect 64 56 65 57 
<< m2 >>
rect 65 56 66 57 
<< m1 >>
rect 66 56 67 57 
<< m2 >>
rect 66 56 67 57 
<< m2c >>
rect 66 56 67 57 
<< m1 >>
rect 66 56 67 57 
<< m2 >>
rect 66 56 67 57 
<< m1 >>
rect 67 56 68 57 
<< m1 >>
rect 70 56 71 57 
<< m2 >>
rect 70 56 71 57 
<< m2c >>
rect 70 56 71 57 
<< m1 >>
rect 70 56 71 57 
<< m2 >>
rect 70 56 71 57 
<< m1 >>
rect 71 56 72 57 
<< m1 >>
rect 72 56 73 57 
<< m1 >>
rect 73 56 74 57 
<< m1 >>
rect 85 56 86 57 
<< m2 >>
rect 85 56 86 57 
<< m2c >>
rect 85 56 86 57 
<< m1 >>
rect 85 56 86 57 
<< m2 >>
rect 85 56 86 57 
<< m1 >>
rect 88 56 89 57 
<< m2 >>
rect 88 56 89 57 
<< m2c >>
rect 88 56 89 57 
<< m1 >>
rect 88 56 89 57 
<< m2 >>
rect 88 56 89 57 
<< m1 >>
rect 89 56 90 57 
<< m1 >>
rect 90 56 91 57 
<< m1 >>
rect 91 56 92 57 
<< m1 >>
rect 98 56 99 57 
<< m2 >>
rect 98 56 99 57 
<< m2c >>
rect 98 56 99 57 
<< m1 >>
rect 98 56 99 57 
<< m2 >>
rect 98 56 99 57 
<< m1 >>
rect 100 56 101 57 
<< m2 >>
rect 100 56 101 57 
<< m2c >>
rect 100 56 101 57 
<< m1 >>
rect 100 56 101 57 
<< m2 >>
rect 100 56 101 57 
<< m2 >>
rect 109 56 110 57 
<< m1 >>
rect 121 56 122 57 
<< m2 >>
rect 121 56 122 57 
<< m2c >>
rect 121 56 122 57 
<< m1 >>
rect 121 56 122 57 
<< m2 >>
rect 121 56 122 57 
<< m1 >>
rect 128 56 129 57 
<< m2 >>
rect 128 56 129 57 
<< m2c >>
rect 128 56 129 57 
<< m1 >>
rect 128 56 129 57 
<< m2 >>
rect 128 56 129 57 
<< m1 >>
rect 136 56 137 57 
<< m1 >>
rect 138 56 139 57 
<< m1 >>
rect 142 56 143 57 
<< m1 >>
rect 145 56 146 57 
<< m1 >>
rect 13 57 14 58 
<< m1 >>
rect 16 57 17 58 
<< m2 >>
rect 30 57 31 58 
<< m2 >>
rect 34 57 35 58 
<< m2 >>
rect 37 57 38 58 
<< m2 >>
rect 52 57 53 58 
<< m2 >>
rect 53 57 54 58 
<< m2 >>
rect 55 57 56 58 
<< m2 >>
rect 57 57 58 58 
<< m1 >>
rect 64 57 65 58 
<< m2 >>
rect 70 57 71 58 
<< m2 >>
rect 85 57 86 58 
<< m2 >>
rect 88 57 89 58 
<< m2 >>
rect 98 57 99 58 
<< m2 >>
rect 100 57 101 58 
<< m2 >>
rect 109 57 110 58 
<< m2 >>
rect 121 57 122 58 
<< m2 >>
rect 128 57 129 58 
<< m1 >>
rect 136 57 137 58 
<< m1 >>
rect 138 57 139 58 
<< m1 >>
rect 142 57 143 58 
<< m1 >>
rect 145 57 146 58 
<< m1 >>
rect 13 58 14 59 
<< m1 >>
rect 16 58 17 59 
<< m1 >>
rect 28 58 29 59 
<< m1 >>
rect 29 58 30 59 
<< m1 >>
rect 30 58 31 59 
<< m2 >>
rect 30 58 31 59 
<< m1 >>
rect 31 58 32 59 
<< m2 >>
rect 31 58 32 59 
<< m1 >>
rect 32 58 33 59 
<< m2 >>
rect 32 58 33 59 
<< m1 >>
rect 33 58 34 59 
<< m2 >>
rect 33 58 34 59 
<< m1 >>
rect 34 58 35 59 
<< m2 >>
rect 34 58 35 59 
<< m1 >>
rect 35 58 36 59 
<< m1 >>
rect 36 58 37 59 
<< m1 >>
rect 37 58 38 59 
<< m2 >>
rect 37 58 38 59 
<< m1 >>
rect 38 58 39 59 
<< m2 >>
rect 38 58 39 59 
<< m1 >>
rect 39 58 40 59 
<< m2 >>
rect 39 58 40 59 
<< m1 >>
rect 40 58 41 59 
<< m2 >>
rect 40 58 41 59 
<< m1 >>
rect 41 58 42 59 
<< m2 >>
rect 41 58 42 59 
<< m1 >>
rect 42 58 43 59 
<< m2 >>
rect 42 58 43 59 
<< m1 >>
rect 43 58 44 59 
<< m2 >>
rect 43 58 44 59 
<< m1 >>
rect 44 58 45 59 
<< m2 >>
rect 44 58 45 59 
<< m1 >>
rect 45 58 46 59 
<< m2 >>
rect 45 58 46 59 
<< m1 >>
rect 46 58 47 59 
<< m2 >>
rect 46 58 47 59 
<< m1 >>
rect 47 58 48 59 
<< m2 >>
rect 47 58 48 59 
<< m1 >>
rect 48 58 49 59 
<< m2 >>
rect 48 58 49 59 
<< m1 >>
rect 49 58 50 59 
<< m2 >>
rect 49 58 50 59 
<< m1 >>
rect 50 58 51 59 
<< m2 >>
rect 50 58 51 59 
<< m1 >>
rect 51 58 52 59 
<< m1 >>
rect 52 58 53 59 
<< m1 >>
rect 53 58 54 59 
<< m2 >>
rect 53 58 54 59 
<< m1 >>
rect 54 58 55 59 
<< m1 >>
rect 55 58 56 59 
<< m2 >>
rect 55 58 56 59 
<< m1 >>
rect 56 58 57 59 
<< m1 >>
rect 57 58 58 59 
<< m2 >>
rect 57 58 58 59 
<< m1 >>
rect 58 58 59 59 
<< m1 >>
rect 59 58 60 59 
<< m1 >>
rect 60 58 61 59 
<< m1 >>
rect 61 58 62 59 
<< m1 >>
rect 62 58 63 59 
<< m2 >>
rect 62 58 63 59 
<< m2c >>
rect 62 58 63 59 
<< m1 >>
rect 62 58 63 59 
<< m2 >>
rect 62 58 63 59 
<< m2 >>
rect 63 58 64 59 
<< m1 >>
rect 64 58 65 59 
<< m2 >>
rect 64 58 65 59 
<< m2 >>
rect 65 58 66 59 
<< m1 >>
rect 66 58 67 59 
<< m2 >>
rect 66 58 67 59 
<< m2c >>
rect 66 58 67 59 
<< m1 >>
rect 66 58 67 59 
<< m2 >>
rect 66 58 67 59 
<< m1 >>
rect 67 58 68 59 
<< m1 >>
rect 68 58 69 59 
<< m1 >>
rect 69 58 70 59 
<< m1 >>
rect 70 58 71 59 
<< m2 >>
rect 70 58 71 59 
<< m1 >>
rect 71 58 72 59 
<< m1 >>
rect 72 58 73 59 
<< m1 >>
rect 73 58 74 59 
<< m1 >>
rect 74 58 75 59 
<< m1 >>
rect 75 58 76 59 
<< m1 >>
rect 76 58 77 59 
<< m1 >>
rect 77 58 78 59 
<< m1 >>
rect 78 58 79 59 
<< m1 >>
rect 79 58 80 59 
<< m1 >>
rect 80 58 81 59 
<< m1 >>
rect 81 58 82 59 
<< m1 >>
rect 82 58 83 59 
<< m1 >>
rect 83 58 84 59 
<< m1 >>
rect 84 58 85 59 
<< m1 >>
rect 85 58 86 59 
<< m2 >>
rect 85 58 86 59 
<< m1 >>
rect 86 58 87 59 
<< m1 >>
rect 87 58 88 59 
<< m1 >>
rect 88 58 89 59 
<< m2 >>
rect 88 58 89 59 
<< m1 >>
rect 89 58 90 59 
<< m1 >>
rect 90 58 91 59 
<< m1 >>
rect 91 58 92 59 
<< m1 >>
rect 92 58 93 59 
<< m1 >>
rect 93 58 94 59 
<< m1 >>
rect 94 58 95 59 
<< m1 >>
rect 95 58 96 59 
<< m1 >>
rect 96 58 97 59 
<< m1 >>
rect 97 58 98 59 
<< m1 >>
rect 98 58 99 59 
<< m2 >>
rect 98 58 99 59 
<< m1 >>
rect 99 58 100 59 
<< m1 >>
rect 100 58 101 59 
<< m2 >>
rect 100 58 101 59 
<< m1 >>
rect 101 58 102 59 
<< m1 >>
rect 102 58 103 59 
<< m1 >>
rect 103 58 104 59 
<< m1 >>
rect 104 58 105 59 
<< m1 >>
rect 105 58 106 59 
<< m1 >>
rect 106 58 107 59 
<< m1 >>
rect 107 58 108 59 
<< m1 >>
rect 108 58 109 59 
<< m1 >>
rect 109 58 110 59 
<< m2 >>
rect 109 58 110 59 
<< m1 >>
rect 110 58 111 59 
<< m1 >>
rect 111 58 112 59 
<< m1 >>
rect 112 58 113 59 
<< m1 >>
rect 113 58 114 59 
<< m1 >>
rect 114 58 115 59 
<< m1 >>
rect 115 58 116 59 
<< m1 >>
rect 116 58 117 59 
<< m1 >>
rect 117 58 118 59 
<< m1 >>
rect 118 58 119 59 
<< m1 >>
rect 119 58 120 59 
<< m1 >>
rect 120 58 121 59 
<< m1 >>
rect 121 58 122 59 
<< m2 >>
rect 121 58 122 59 
<< m1 >>
rect 122 58 123 59 
<< m1 >>
rect 123 58 124 59 
<< m1 >>
rect 124 58 125 59 
<< m1 >>
rect 125 58 126 59 
<< m1 >>
rect 126 58 127 59 
<< m1 >>
rect 127 58 128 59 
<< m1 >>
rect 128 58 129 59 
<< m2 >>
rect 128 58 129 59 
<< m1 >>
rect 129 58 130 59 
<< m1 >>
rect 130 58 131 59 
<< m1 >>
rect 131 58 132 59 
<< m1 >>
rect 132 58 133 59 
<< m1 >>
rect 133 58 134 59 
<< m1 >>
rect 134 58 135 59 
<< m1 >>
rect 135 58 136 59 
<< m1 >>
rect 136 58 137 59 
<< m1 >>
rect 138 58 139 59 
<< m1 >>
rect 139 58 140 59 
<< m1 >>
rect 140 58 141 59 
<< m1 >>
rect 141 58 142 59 
<< m1 >>
rect 142 58 143 59 
<< m1 >>
rect 145 58 146 59 
<< m1 >>
rect 13 59 14 60 
<< m1 >>
rect 16 59 17 60 
<< m1 >>
rect 28 59 29 60 
<< m2 >>
rect 50 59 51 60 
<< m2 >>
rect 53 59 54 60 
<< m2 >>
rect 55 59 56 60 
<< m2 >>
rect 57 59 58 60 
<< m1 >>
rect 64 59 65 60 
<< m2 >>
rect 70 59 71 60 
<< m2 >>
rect 85 59 86 60 
<< m2 >>
rect 88 59 89 60 
<< m2 >>
rect 98 59 99 60 
<< m2 >>
rect 100 59 101 60 
<< m2 >>
rect 109 59 110 60 
<< m2 >>
rect 121 59 122 60 
<< m2 >>
rect 128 59 129 60 
<< m1 >>
rect 145 59 146 60 
<< m1 >>
rect 13 60 14 61 
<< m1 >>
rect 16 60 17 61 
<< m1 >>
rect 17 60 18 61 
<< m1 >>
rect 18 60 19 61 
<< m1 >>
rect 19 60 20 61 
<< m1 >>
rect 20 60 21 61 
<< m1 >>
rect 21 60 22 61 
<< m1 >>
rect 22 60 23 61 
<< m1 >>
rect 23 60 24 61 
<< m1 >>
rect 24 60 25 61 
<< m1 >>
rect 25 60 26 61 
<< m1 >>
rect 26 60 27 61 
<< m2 >>
rect 26 60 27 61 
<< m2c >>
rect 26 60 27 61 
<< m1 >>
rect 26 60 27 61 
<< m2 >>
rect 26 60 27 61 
<< m2 >>
rect 27 60 28 61 
<< m1 >>
rect 28 60 29 61 
<< m2 >>
rect 28 60 29 61 
<< m2 >>
rect 29 60 30 61 
<< m1 >>
rect 30 60 31 61 
<< m2 >>
rect 30 60 31 61 
<< m2c >>
rect 30 60 31 61 
<< m1 >>
rect 30 60 31 61 
<< m2 >>
rect 30 60 31 61 
<< m1 >>
rect 31 60 32 61 
<< m1 >>
rect 32 60 33 61 
<< m1 >>
rect 33 60 34 61 
<< m1 >>
rect 34 60 35 61 
<< m1 >>
rect 35 60 36 61 
<< m1 >>
rect 36 60 37 61 
<< m1 >>
rect 37 60 38 61 
<< m1 >>
rect 38 60 39 61 
<< m1 >>
rect 39 60 40 61 
<< m1 >>
rect 40 60 41 61 
<< m1 >>
rect 41 60 42 61 
<< m1 >>
rect 42 60 43 61 
<< m1 >>
rect 43 60 44 61 
<< m1 >>
rect 44 60 45 61 
<< m1 >>
rect 45 60 46 61 
<< m1 >>
rect 46 60 47 61 
<< m1 >>
rect 47 60 48 61 
<< m1 >>
rect 48 60 49 61 
<< m1 >>
rect 49 60 50 61 
<< m1 >>
rect 50 60 51 61 
<< m2 >>
rect 50 60 51 61 
<< m1 >>
rect 51 60 52 61 
<< m1 >>
rect 52 60 53 61 
<< m1 >>
rect 53 60 54 61 
<< m2 >>
rect 53 60 54 61 
<< m1 >>
rect 54 60 55 61 
<< m1 >>
rect 55 60 56 61 
<< m2 >>
rect 55 60 56 61 
<< m1 >>
rect 56 60 57 61 
<< m1 >>
rect 57 60 58 61 
<< m2 >>
rect 57 60 58 61 
<< m1 >>
rect 58 60 59 61 
<< m1 >>
rect 59 60 60 61 
<< m1 >>
rect 60 60 61 61 
<< m1 >>
rect 61 60 62 61 
<< m1 >>
rect 62 60 63 61 
<< m2 >>
rect 62 60 63 61 
<< m2c >>
rect 62 60 63 61 
<< m1 >>
rect 62 60 63 61 
<< m2 >>
rect 62 60 63 61 
<< m2 >>
rect 63 60 64 61 
<< m1 >>
rect 64 60 65 61 
<< m2 >>
rect 64 60 65 61 
<< m2 >>
rect 65 60 66 61 
<< m1 >>
rect 66 60 67 61 
<< m2 >>
rect 66 60 67 61 
<< m2c >>
rect 66 60 67 61 
<< m1 >>
rect 66 60 67 61 
<< m2 >>
rect 66 60 67 61 
<< m1 >>
rect 67 60 68 61 
<< m1 >>
rect 68 60 69 61 
<< m1 >>
rect 69 60 70 61 
<< m1 >>
rect 70 60 71 61 
<< m2 >>
rect 70 60 71 61 
<< m1 >>
rect 71 60 72 61 
<< m1 >>
rect 72 60 73 61 
<< m1 >>
rect 73 60 74 61 
<< m1 >>
rect 74 60 75 61 
<< m1 >>
rect 75 60 76 61 
<< m1 >>
rect 76 60 77 61 
<< m1 >>
rect 77 60 78 61 
<< m1 >>
rect 78 60 79 61 
<< m1 >>
rect 79 60 80 61 
<< m1 >>
rect 80 60 81 61 
<< m1 >>
rect 81 60 82 61 
<< m1 >>
rect 82 60 83 61 
<< m1 >>
rect 83 60 84 61 
<< m1 >>
rect 84 60 85 61 
<< m1 >>
rect 85 60 86 61 
<< m2 >>
rect 85 60 86 61 
<< m2c >>
rect 85 60 86 61 
<< m1 >>
rect 85 60 86 61 
<< m2 >>
rect 85 60 86 61 
<< m1 >>
rect 88 60 89 61 
<< m2 >>
rect 88 60 89 61 
<< m2c >>
rect 88 60 89 61 
<< m1 >>
rect 88 60 89 61 
<< m2 >>
rect 88 60 89 61 
<< m1 >>
rect 98 60 99 61 
<< m2 >>
rect 98 60 99 61 
<< m2c >>
rect 98 60 99 61 
<< m1 >>
rect 98 60 99 61 
<< m2 >>
rect 98 60 99 61 
<< m1 >>
rect 100 60 101 61 
<< m2 >>
rect 100 60 101 61 
<< m2c >>
rect 100 60 101 61 
<< m1 >>
rect 100 60 101 61 
<< m2 >>
rect 100 60 101 61 
<< m1 >>
rect 106 60 107 61 
<< m1 >>
rect 107 60 108 61 
<< m1 >>
rect 108 60 109 61 
<< m1 >>
rect 109 60 110 61 
<< m2 >>
rect 109 60 110 61 
<< m1 >>
rect 110 60 111 61 
<< m1 >>
rect 111 60 112 61 
<< m1 >>
rect 112 60 113 61 
<< m1 >>
rect 113 60 114 61 
<< m1 >>
rect 114 60 115 61 
<< m1 >>
rect 115 60 116 61 
<< m1 >>
rect 116 60 117 61 
<< m1 >>
rect 117 60 118 61 
<< m1 >>
rect 118 60 119 61 
<< m1 >>
rect 119 60 120 61 
<< m1 >>
rect 120 60 121 61 
<< m1 >>
rect 121 60 122 61 
<< m2 >>
rect 121 60 122 61 
<< m2c >>
rect 121 60 122 61 
<< m1 >>
rect 121 60 122 61 
<< m2 >>
rect 121 60 122 61 
<< m1 >>
rect 128 60 129 61 
<< m2 >>
rect 128 60 129 61 
<< m2c >>
rect 128 60 129 61 
<< m1 >>
rect 128 60 129 61 
<< m2 >>
rect 128 60 129 61 
<< m1 >>
rect 129 60 130 61 
<< m1 >>
rect 145 60 146 61 
<< m1 >>
rect 10 61 11 62 
<< m1 >>
rect 11 61 12 62 
<< m1 >>
rect 12 61 13 62 
<< m1 >>
rect 13 61 14 62 
<< m1 >>
rect 28 61 29 62 
<< m2 >>
rect 50 61 51 62 
<< m2 >>
rect 53 61 54 62 
<< m2 >>
rect 55 61 56 62 
<< m2 >>
rect 57 61 58 62 
<< m1 >>
rect 64 61 65 62 
<< m2 >>
rect 70 61 71 62 
<< m1 >>
rect 88 61 89 62 
<< m1 >>
rect 98 61 99 62 
<< m1 >>
rect 100 61 101 62 
<< m1 >>
rect 102 61 103 62 
<< m1 >>
rect 103 61 104 62 
<< m1 >>
rect 104 61 105 62 
<< m2 >>
rect 104 61 105 62 
<< m2c >>
rect 104 61 105 62 
<< m1 >>
rect 104 61 105 62 
<< m2 >>
rect 104 61 105 62 
<< m2 >>
rect 105 61 106 62 
<< m1 >>
rect 106 61 107 62 
<< m2 >>
rect 106 61 107 62 
<< m2 >>
rect 107 61 108 62 
<< m2 >>
rect 108 61 109 62 
<< m2 >>
rect 109 61 110 62 
<< m1 >>
rect 129 61 130 62 
<< m1 >>
rect 145 61 146 62 
<< m1 >>
rect 10 62 11 63 
<< m1 >>
rect 28 62 29 63 
<< m1 >>
rect 50 62 51 63 
<< m2 >>
rect 50 62 51 63 
<< m2c >>
rect 50 62 51 63 
<< m1 >>
rect 50 62 51 63 
<< m2 >>
rect 50 62 51 63 
<< m1 >>
rect 51 62 52 63 
<< m1 >>
rect 52 62 53 63 
<< m1 >>
rect 53 62 54 63 
<< m2 >>
rect 53 62 54 63 
<< m1 >>
rect 54 62 55 63 
<< m1 >>
rect 55 62 56 63 
<< m2 >>
rect 55 62 56 63 
<< m1 >>
rect 56 62 57 63 
<< m1 >>
rect 57 62 58 63 
<< m2 >>
rect 57 62 58 63 
<< m1 >>
rect 58 62 59 63 
<< m1 >>
rect 59 62 60 63 
<< m1 >>
rect 60 62 61 63 
<< m1 >>
rect 61 62 62 63 
<< m1 >>
rect 62 62 63 63 
<< m2 >>
rect 62 62 63 63 
<< m2c >>
rect 62 62 63 63 
<< m1 >>
rect 62 62 63 63 
<< m2 >>
rect 62 62 63 63 
<< m2 >>
rect 63 62 64 63 
<< m1 >>
rect 64 62 65 63 
<< m1 >>
rect 70 62 71 63 
<< m2 >>
rect 70 62 71 63 
<< m2c >>
rect 70 62 71 63 
<< m1 >>
rect 70 62 71 63 
<< m2 >>
rect 70 62 71 63 
<< m1 >>
rect 88 62 89 63 
<< m1 >>
rect 98 62 99 63 
<< m1 >>
rect 100 62 101 63 
<< m1 >>
rect 102 62 103 63 
<< m1 >>
rect 106 62 107 63 
<< m1 >>
rect 129 62 130 63 
<< m1 >>
rect 145 62 146 63 
<< m1 >>
rect 10 63 11 64 
<< m1 >>
rect 28 63 29 64 
<< m2 >>
rect 53 63 54 64 
<< m2 >>
rect 55 63 56 64 
<< m2 >>
rect 57 63 58 64 
<< m2 >>
rect 63 63 64 64 
<< m1 >>
rect 64 63 65 64 
<< m1 >>
rect 70 63 71 64 
<< m2 >>
rect 87 63 88 64 
<< m1 >>
rect 88 63 89 64 
<< m2 >>
rect 88 63 89 64 
<< m2 >>
rect 89 63 90 64 
<< m1 >>
rect 90 63 91 64 
<< m2 >>
rect 90 63 91 64 
<< m2c >>
rect 90 63 91 64 
<< m1 >>
rect 90 63 91 64 
<< m2 >>
rect 90 63 91 64 
<< m1 >>
rect 91 63 92 64 
<< m1 >>
rect 92 63 93 64 
<< m1 >>
rect 93 63 94 64 
<< m1 >>
rect 94 63 95 64 
<< m1 >>
rect 95 63 96 64 
<< m1 >>
rect 96 63 97 64 
<< m2 >>
rect 96 63 97 64 
<< m2c >>
rect 96 63 97 64 
<< m1 >>
rect 96 63 97 64 
<< m2 >>
rect 96 63 97 64 
<< m2 >>
rect 97 63 98 64 
<< m1 >>
rect 98 63 99 64 
<< m2 >>
rect 98 63 99 64 
<< m2 >>
rect 99 63 100 64 
<< m1 >>
rect 100 63 101 64 
<< m2 >>
rect 100 63 101 64 
<< m2 >>
rect 101 63 102 64 
<< m1 >>
rect 102 63 103 64 
<< m2 >>
rect 102 63 103 64 
<< m2c >>
rect 102 63 103 64 
<< m1 >>
rect 102 63 103 64 
<< m2 >>
rect 102 63 103 64 
<< m1 >>
rect 106 63 107 64 
<< m1 >>
rect 129 63 130 64 
<< m1 >>
rect 145 63 146 64 
<< m1 >>
rect 10 64 11 65 
<< m1 >>
rect 24 64 25 65 
<< m1 >>
rect 25 64 26 65 
<< m1 >>
rect 26 64 27 65 
<< m2 >>
rect 26 64 27 65 
<< m2c >>
rect 26 64 27 65 
<< m1 >>
rect 26 64 27 65 
<< m2 >>
rect 26 64 27 65 
<< m2 >>
rect 27 64 28 65 
<< m1 >>
rect 28 64 29 65 
<< m2 >>
rect 28 64 29 65 
<< m2 >>
rect 29 64 30 65 
<< m1 >>
rect 30 64 31 65 
<< m2 >>
rect 30 64 31 65 
<< m2c >>
rect 30 64 31 65 
<< m1 >>
rect 30 64 31 65 
<< m2 >>
rect 30 64 31 65 
<< m1 >>
rect 31 64 32 65 
<< m1 >>
rect 53 64 54 65 
<< m2 >>
rect 53 64 54 65 
<< m2c >>
rect 53 64 54 65 
<< m1 >>
rect 53 64 54 65 
<< m2 >>
rect 53 64 54 65 
<< m1 >>
rect 54 64 55 65 
<< m1 >>
rect 55 64 56 65 
<< m2 >>
rect 55 64 56 65 
<< m1 >>
rect 57 64 58 65 
<< m2 >>
rect 57 64 58 65 
<< m2c >>
rect 57 64 58 65 
<< m1 >>
rect 57 64 58 65 
<< m2 >>
rect 57 64 58 65 
<< m2 >>
rect 63 64 64 65 
<< m1 >>
rect 64 64 65 65 
<< m1 >>
rect 70 64 71 65 
<< m1 >>
rect 85 64 86 65 
<< m1 >>
rect 86 64 87 65 
<< m2 >>
rect 86 64 87 65 
<< m2c >>
rect 86 64 87 65 
<< m1 >>
rect 86 64 87 65 
<< m2 >>
rect 86 64 87 65 
<< m2 >>
rect 87 64 88 65 
<< m1 >>
rect 88 64 89 65 
<< m1 >>
rect 98 64 99 65 
<< m1 >>
rect 100 64 101 65 
<< m1 >>
rect 106 64 107 65 
<< m1 >>
rect 118 64 119 65 
<< m1 >>
rect 119 64 120 65 
<< m1 >>
rect 120 64 121 65 
<< m1 >>
rect 121 64 122 65 
<< m1 >>
rect 124 64 125 65 
<< m1 >>
rect 125 64 126 65 
<< m1 >>
rect 126 64 127 65 
<< m1 >>
rect 127 64 128 65 
<< m1 >>
rect 129 64 130 65 
<< m1 >>
rect 145 64 146 65 
<< m1 >>
rect 10 65 11 66 
<< m1 >>
rect 24 65 25 66 
<< m1 >>
rect 28 65 29 66 
<< m1 >>
rect 31 65 32 66 
<< m1 >>
rect 55 65 56 66 
<< m2 >>
rect 55 65 56 66 
<< m1 >>
rect 57 65 58 66 
<< m2 >>
rect 63 65 64 66 
<< m1 >>
rect 64 65 65 66 
<< m1 >>
rect 70 65 71 66 
<< m1 >>
rect 85 65 86 66 
<< m1 >>
rect 88 65 89 66 
<< m1 >>
rect 98 65 99 66 
<< m1 >>
rect 100 65 101 66 
<< m1 >>
rect 106 65 107 66 
<< m1 >>
rect 118 65 119 66 
<< m1 >>
rect 121 65 122 66 
<< m1 >>
rect 124 65 125 66 
<< m1 >>
rect 127 65 128 66 
<< m1 >>
rect 129 65 130 66 
<< m1 >>
rect 145 65 146 66 
<< m1 >>
rect 10 66 11 67 
<< pdiffusion >>
rect 12 66 13 67 
<< pdiffusion >>
rect 13 66 14 67 
<< pdiffusion >>
rect 14 66 15 67 
<< pdiffusion >>
rect 15 66 16 67 
<< pdiffusion >>
rect 16 66 17 67 
<< pdiffusion >>
rect 17 66 18 67 
<< m1 >>
rect 24 66 25 67 
<< m1 >>
rect 28 66 29 67 
<< pdiffusion >>
rect 30 66 31 67 
<< m1 >>
rect 31 66 32 67 
<< pdiffusion >>
rect 31 66 32 67 
<< pdiffusion >>
rect 32 66 33 67 
<< pdiffusion >>
rect 33 66 34 67 
<< pdiffusion >>
rect 34 66 35 67 
<< pdiffusion >>
rect 35 66 36 67 
<< pdiffusion >>
rect 48 66 49 67 
<< pdiffusion >>
rect 49 66 50 67 
<< pdiffusion >>
rect 50 66 51 67 
<< pdiffusion >>
rect 51 66 52 67 
<< pdiffusion >>
rect 52 66 53 67 
<< pdiffusion >>
rect 53 66 54 67 
<< m1 >>
rect 55 66 56 67 
<< m2 >>
rect 55 66 56 67 
<< m1 >>
rect 57 66 58 67 
<< m2 >>
rect 63 66 64 67 
<< m1 >>
rect 64 66 65 67 
<< pdiffusion >>
rect 66 66 67 67 
<< pdiffusion >>
rect 67 66 68 67 
<< pdiffusion >>
rect 68 66 69 67 
<< pdiffusion >>
rect 69 66 70 67 
<< m1 >>
rect 70 66 71 67 
<< pdiffusion >>
rect 70 66 71 67 
<< pdiffusion >>
rect 71 66 72 67 
<< pdiffusion >>
rect 84 66 85 67 
<< m1 >>
rect 85 66 86 67 
<< pdiffusion >>
rect 85 66 86 67 
<< pdiffusion >>
rect 86 66 87 67 
<< pdiffusion >>
rect 87 66 88 67 
<< m1 >>
rect 88 66 89 67 
<< pdiffusion >>
rect 88 66 89 67 
<< pdiffusion >>
rect 89 66 90 67 
<< m1 >>
rect 98 66 99 67 
<< m1 >>
rect 100 66 101 67 
<< pdiffusion >>
rect 102 66 103 67 
<< pdiffusion >>
rect 103 66 104 67 
<< pdiffusion >>
rect 104 66 105 67 
<< pdiffusion >>
rect 105 66 106 67 
<< m1 >>
rect 106 66 107 67 
<< pdiffusion >>
rect 106 66 107 67 
<< pdiffusion >>
rect 107 66 108 67 
<< m1 >>
rect 118 66 119 67 
<< pdiffusion >>
rect 120 66 121 67 
<< m1 >>
rect 121 66 122 67 
<< pdiffusion >>
rect 121 66 122 67 
<< pdiffusion >>
rect 122 66 123 67 
<< pdiffusion >>
rect 123 66 124 67 
<< m1 >>
rect 124 66 125 67 
<< pdiffusion >>
rect 124 66 125 67 
<< pdiffusion >>
rect 125 66 126 67 
<< m1 >>
rect 127 66 128 67 
<< m1 >>
rect 129 66 130 67 
<< pdiffusion >>
rect 138 66 139 67 
<< pdiffusion >>
rect 139 66 140 67 
<< pdiffusion >>
rect 140 66 141 67 
<< pdiffusion >>
rect 141 66 142 67 
<< pdiffusion >>
rect 142 66 143 67 
<< pdiffusion >>
rect 143 66 144 67 
<< m1 >>
rect 145 66 146 67 
<< m1 >>
rect 10 67 11 68 
<< pdiffusion >>
rect 12 67 13 68 
<< pdiffusion >>
rect 13 67 14 68 
<< pdiffusion >>
rect 14 67 15 68 
<< pdiffusion >>
rect 15 67 16 68 
<< pdiffusion >>
rect 16 67 17 68 
<< pdiffusion >>
rect 17 67 18 68 
<< m1 >>
rect 24 67 25 68 
<< m1 >>
rect 28 67 29 68 
<< pdiffusion >>
rect 30 67 31 68 
<< pdiffusion >>
rect 31 67 32 68 
<< pdiffusion >>
rect 32 67 33 68 
<< pdiffusion >>
rect 33 67 34 68 
<< pdiffusion >>
rect 34 67 35 68 
<< pdiffusion >>
rect 35 67 36 68 
<< pdiffusion >>
rect 48 67 49 68 
<< pdiffusion >>
rect 49 67 50 68 
<< pdiffusion >>
rect 50 67 51 68 
<< pdiffusion >>
rect 51 67 52 68 
<< pdiffusion >>
rect 52 67 53 68 
<< pdiffusion >>
rect 53 67 54 68 
<< m1 >>
rect 55 67 56 68 
<< m2 >>
rect 55 67 56 68 
<< m1 >>
rect 57 67 58 68 
<< m2 >>
rect 63 67 64 68 
<< m1 >>
rect 64 67 65 68 
<< pdiffusion >>
rect 66 67 67 68 
<< pdiffusion >>
rect 67 67 68 68 
<< pdiffusion >>
rect 68 67 69 68 
<< pdiffusion >>
rect 69 67 70 68 
<< pdiffusion >>
rect 70 67 71 68 
<< pdiffusion >>
rect 71 67 72 68 
<< pdiffusion >>
rect 84 67 85 68 
<< pdiffusion >>
rect 85 67 86 68 
<< pdiffusion >>
rect 86 67 87 68 
<< pdiffusion >>
rect 87 67 88 68 
<< pdiffusion >>
rect 88 67 89 68 
<< pdiffusion >>
rect 89 67 90 68 
<< m1 >>
rect 98 67 99 68 
<< m1 >>
rect 100 67 101 68 
<< pdiffusion >>
rect 102 67 103 68 
<< pdiffusion >>
rect 103 67 104 68 
<< pdiffusion >>
rect 104 67 105 68 
<< pdiffusion >>
rect 105 67 106 68 
<< pdiffusion >>
rect 106 67 107 68 
<< pdiffusion >>
rect 107 67 108 68 
<< m1 >>
rect 118 67 119 68 
<< pdiffusion >>
rect 120 67 121 68 
<< pdiffusion >>
rect 121 67 122 68 
<< pdiffusion >>
rect 122 67 123 68 
<< pdiffusion >>
rect 123 67 124 68 
<< pdiffusion >>
rect 124 67 125 68 
<< pdiffusion >>
rect 125 67 126 68 
<< m1 >>
rect 127 67 128 68 
<< m1 >>
rect 129 67 130 68 
<< pdiffusion >>
rect 138 67 139 68 
<< pdiffusion >>
rect 139 67 140 68 
<< pdiffusion >>
rect 140 67 141 68 
<< pdiffusion >>
rect 141 67 142 68 
<< pdiffusion >>
rect 142 67 143 68 
<< pdiffusion >>
rect 143 67 144 68 
<< m1 >>
rect 145 67 146 68 
<< m1 >>
rect 10 68 11 69 
<< pdiffusion >>
rect 12 68 13 69 
<< pdiffusion >>
rect 13 68 14 69 
<< pdiffusion >>
rect 14 68 15 69 
<< pdiffusion >>
rect 15 68 16 69 
<< pdiffusion >>
rect 16 68 17 69 
<< pdiffusion >>
rect 17 68 18 69 
<< m1 >>
rect 24 68 25 69 
<< m1 >>
rect 28 68 29 69 
<< pdiffusion >>
rect 30 68 31 69 
<< pdiffusion >>
rect 31 68 32 69 
<< pdiffusion >>
rect 32 68 33 69 
<< pdiffusion >>
rect 33 68 34 69 
<< pdiffusion >>
rect 34 68 35 69 
<< pdiffusion >>
rect 35 68 36 69 
<< pdiffusion >>
rect 48 68 49 69 
<< pdiffusion >>
rect 49 68 50 69 
<< pdiffusion >>
rect 50 68 51 69 
<< pdiffusion >>
rect 51 68 52 69 
<< pdiffusion >>
rect 52 68 53 69 
<< pdiffusion >>
rect 53 68 54 69 
<< m1 >>
rect 55 68 56 69 
<< m2 >>
rect 55 68 56 69 
<< m1 >>
rect 57 68 58 69 
<< m2 >>
rect 63 68 64 69 
<< m1 >>
rect 64 68 65 69 
<< pdiffusion >>
rect 66 68 67 69 
<< pdiffusion >>
rect 67 68 68 69 
<< pdiffusion >>
rect 68 68 69 69 
<< pdiffusion >>
rect 69 68 70 69 
<< pdiffusion >>
rect 70 68 71 69 
<< pdiffusion >>
rect 71 68 72 69 
<< pdiffusion >>
rect 84 68 85 69 
<< pdiffusion >>
rect 85 68 86 69 
<< pdiffusion >>
rect 86 68 87 69 
<< pdiffusion >>
rect 87 68 88 69 
<< pdiffusion >>
rect 88 68 89 69 
<< pdiffusion >>
rect 89 68 90 69 
<< m1 >>
rect 98 68 99 69 
<< m1 >>
rect 100 68 101 69 
<< pdiffusion >>
rect 102 68 103 69 
<< pdiffusion >>
rect 103 68 104 69 
<< pdiffusion >>
rect 104 68 105 69 
<< pdiffusion >>
rect 105 68 106 69 
<< pdiffusion >>
rect 106 68 107 69 
<< pdiffusion >>
rect 107 68 108 69 
<< m1 >>
rect 118 68 119 69 
<< pdiffusion >>
rect 120 68 121 69 
<< pdiffusion >>
rect 121 68 122 69 
<< pdiffusion >>
rect 122 68 123 69 
<< pdiffusion >>
rect 123 68 124 69 
<< pdiffusion >>
rect 124 68 125 69 
<< pdiffusion >>
rect 125 68 126 69 
<< m1 >>
rect 127 68 128 69 
<< m1 >>
rect 129 68 130 69 
<< pdiffusion >>
rect 138 68 139 69 
<< pdiffusion >>
rect 139 68 140 69 
<< pdiffusion >>
rect 140 68 141 69 
<< pdiffusion >>
rect 141 68 142 69 
<< pdiffusion >>
rect 142 68 143 69 
<< pdiffusion >>
rect 143 68 144 69 
<< m1 >>
rect 145 68 146 69 
<< m1 >>
rect 10 69 11 70 
<< pdiffusion >>
rect 12 69 13 70 
<< pdiffusion >>
rect 13 69 14 70 
<< pdiffusion >>
rect 14 69 15 70 
<< pdiffusion >>
rect 15 69 16 70 
<< pdiffusion >>
rect 16 69 17 70 
<< pdiffusion >>
rect 17 69 18 70 
<< m1 >>
rect 24 69 25 70 
<< m1 >>
rect 28 69 29 70 
<< pdiffusion >>
rect 30 69 31 70 
<< pdiffusion >>
rect 31 69 32 70 
<< pdiffusion >>
rect 32 69 33 70 
<< pdiffusion >>
rect 33 69 34 70 
<< pdiffusion >>
rect 34 69 35 70 
<< pdiffusion >>
rect 35 69 36 70 
<< pdiffusion >>
rect 48 69 49 70 
<< pdiffusion >>
rect 49 69 50 70 
<< pdiffusion >>
rect 50 69 51 70 
<< pdiffusion >>
rect 51 69 52 70 
<< pdiffusion >>
rect 52 69 53 70 
<< pdiffusion >>
rect 53 69 54 70 
<< m1 >>
rect 55 69 56 70 
<< m2 >>
rect 55 69 56 70 
<< m1 >>
rect 57 69 58 70 
<< m2 >>
rect 63 69 64 70 
<< m1 >>
rect 64 69 65 70 
<< pdiffusion >>
rect 66 69 67 70 
<< pdiffusion >>
rect 67 69 68 70 
<< pdiffusion >>
rect 68 69 69 70 
<< pdiffusion >>
rect 69 69 70 70 
<< pdiffusion >>
rect 70 69 71 70 
<< pdiffusion >>
rect 71 69 72 70 
<< pdiffusion >>
rect 84 69 85 70 
<< pdiffusion >>
rect 85 69 86 70 
<< pdiffusion >>
rect 86 69 87 70 
<< pdiffusion >>
rect 87 69 88 70 
<< pdiffusion >>
rect 88 69 89 70 
<< pdiffusion >>
rect 89 69 90 70 
<< m1 >>
rect 98 69 99 70 
<< m1 >>
rect 100 69 101 70 
<< pdiffusion >>
rect 102 69 103 70 
<< pdiffusion >>
rect 103 69 104 70 
<< pdiffusion >>
rect 104 69 105 70 
<< pdiffusion >>
rect 105 69 106 70 
<< pdiffusion >>
rect 106 69 107 70 
<< pdiffusion >>
rect 107 69 108 70 
<< m1 >>
rect 118 69 119 70 
<< pdiffusion >>
rect 120 69 121 70 
<< pdiffusion >>
rect 121 69 122 70 
<< pdiffusion >>
rect 122 69 123 70 
<< pdiffusion >>
rect 123 69 124 70 
<< pdiffusion >>
rect 124 69 125 70 
<< pdiffusion >>
rect 125 69 126 70 
<< m1 >>
rect 127 69 128 70 
<< m1 >>
rect 129 69 130 70 
<< pdiffusion >>
rect 138 69 139 70 
<< pdiffusion >>
rect 139 69 140 70 
<< pdiffusion >>
rect 140 69 141 70 
<< pdiffusion >>
rect 141 69 142 70 
<< pdiffusion >>
rect 142 69 143 70 
<< pdiffusion >>
rect 143 69 144 70 
<< m1 >>
rect 145 69 146 70 
<< m1 >>
rect 10 70 11 71 
<< pdiffusion >>
rect 12 70 13 71 
<< pdiffusion >>
rect 13 70 14 71 
<< pdiffusion >>
rect 14 70 15 71 
<< pdiffusion >>
rect 15 70 16 71 
<< pdiffusion >>
rect 16 70 17 71 
<< pdiffusion >>
rect 17 70 18 71 
<< m1 >>
rect 24 70 25 71 
<< m1 >>
rect 28 70 29 71 
<< pdiffusion >>
rect 30 70 31 71 
<< pdiffusion >>
rect 31 70 32 71 
<< pdiffusion >>
rect 32 70 33 71 
<< pdiffusion >>
rect 33 70 34 71 
<< pdiffusion >>
rect 34 70 35 71 
<< pdiffusion >>
rect 35 70 36 71 
<< pdiffusion >>
rect 48 70 49 71 
<< pdiffusion >>
rect 49 70 50 71 
<< pdiffusion >>
rect 50 70 51 71 
<< pdiffusion >>
rect 51 70 52 71 
<< pdiffusion >>
rect 52 70 53 71 
<< pdiffusion >>
rect 53 70 54 71 
<< m1 >>
rect 55 70 56 71 
<< m2 >>
rect 55 70 56 71 
<< m1 >>
rect 57 70 58 71 
<< m2 >>
rect 63 70 64 71 
<< m1 >>
rect 64 70 65 71 
<< pdiffusion >>
rect 66 70 67 71 
<< pdiffusion >>
rect 67 70 68 71 
<< pdiffusion >>
rect 68 70 69 71 
<< pdiffusion >>
rect 69 70 70 71 
<< pdiffusion >>
rect 70 70 71 71 
<< pdiffusion >>
rect 71 70 72 71 
<< pdiffusion >>
rect 84 70 85 71 
<< pdiffusion >>
rect 85 70 86 71 
<< pdiffusion >>
rect 86 70 87 71 
<< pdiffusion >>
rect 87 70 88 71 
<< pdiffusion >>
rect 88 70 89 71 
<< pdiffusion >>
rect 89 70 90 71 
<< m1 >>
rect 98 70 99 71 
<< m1 >>
rect 100 70 101 71 
<< pdiffusion >>
rect 102 70 103 71 
<< pdiffusion >>
rect 103 70 104 71 
<< pdiffusion >>
rect 104 70 105 71 
<< pdiffusion >>
rect 105 70 106 71 
<< pdiffusion >>
rect 106 70 107 71 
<< pdiffusion >>
rect 107 70 108 71 
<< m1 >>
rect 118 70 119 71 
<< pdiffusion >>
rect 120 70 121 71 
<< pdiffusion >>
rect 121 70 122 71 
<< pdiffusion >>
rect 122 70 123 71 
<< pdiffusion >>
rect 123 70 124 71 
<< pdiffusion >>
rect 124 70 125 71 
<< pdiffusion >>
rect 125 70 126 71 
<< m1 >>
rect 127 70 128 71 
<< m1 >>
rect 129 70 130 71 
<< pdiffusion >>
rect 138 70 139 71 
<< pdiffusion >>
rect 139 70 140 71 
<< pdiffusion >>
rect 140 70 141 71 
<< pdiffusion >>
rect 141 70 142 71 
<< pdiffusion >>
rect 142 70 143 71 
<< pdiffusion >>
rect 143 70 144 71 
<< m1 >>
rect 145 70 146 71 
<< m1 >>
rect 10 71 11 72 
<< pdiffusion >>
rect 12 71 13 72 
<< m1 >>
rect 13 71 14 72 
<< pdiffusion >>
rect 13 71 14 72 
<< pdiffusion >>
rect 14 71 15 72 
<< pdiffusion >>
rect 15 71 16 72 
<< m1 >>
rect 16 71 17 72 
<< pdiffusion >>
rect 16 71 17 72 
<< pdiffusion >>
rect 17 71 18 72 
<< m1 >>
rect 24 71 25 72 
<< m2 >>
rect 24 71 25 72 
<< m2c >>
rect 24 71 25 72 
<< m1 >>
rect 24 71 25 72 
<< m2 >>
rect 24 71 25 72 
<< m1 >>
rect 28 71 29 72 
<< pdiffusion >>
rect 30 71 31 72 
<< pdiffusion >>
rect 31 71 32 72 
<< pdiffusion >>
rect 32 71 33 72 
<< pdiffusion >>
rect 33 71 34 72 
<< m1 >>
rect 34 71 35 72 
<< pdiffusion >>
rect 34 71 35 72 
<< pdiffusion >>
rect 35 71 36 72 
<< pdiffusion >>
rect 48 71 49 72 
<< m1 >>
rect 49 71 50 72 
<< pdiffusion >>
rect 49 71 50 72 
<< pdiffusion >>
rect 50 71 51 72 
<< pdiffusion >>
rect 51 71 52 72 
<< m1 >>
rect 52 71 53 72 
<< pdiffusion >>
rect 52 71 53 72 
<< pdiffusion >>
rect 53 71 54 72 
<< m1 >>
rect 55 71 56 72 
<< m2 >>
rect 55 71 56 72 
<< m1 >>
rect 57 71 58 72 
<< m2 >>
rect 63 71 64 72 
<< m1 >>
rect 64 71 65 72 
<< pdiffusion >>
rect 66 71 67 72 
<< pdiffusion >>
rect 67 71 68 72 
<< pdiffusion >>
rect 68 71 69 72 
<< pdiffusion >>
rect 69 71 70 72 
<< pdiffusion >>
rect 70 71 71 72 
<< pdiffusion >>
rect 71 71 72 72 
<< pdiffusion >>
rect 84 71 85 72 
<< pdiffusion >>
rect 85 71 86 72 
<< pdiffusion >>
rect 86 71 87 72 
<< pdiffusion >>
rect 87 71 88 72 
<< m1 >>
rect 88 71 89 72 
<< pdiffusion >>
rect 88 71 89 72 
<< pdiffusion >>
rect 89 71 90 72 
<< m1 >>
rect 98 71 99 72 
<< m1 >>
rect 100 71 101 72 
<< pdiffusion >>
rect 102 71 103 72 
<< m1 >>
rect 103 71 104 72 
<< pdiffusion >>
rect 103 71 104 72 
<< pdiffusion >>
rect 104 71 105 72 
<< pdiffusion >>
rect 105 71 106 72 
<< pdiffusion >>
rect 106 71 107 72 
<< pdiffusion >>
rect 107 71 108 72 
<< m1 >>
rect 118 71 119 72 
<< pdiffusion >>
rect 120 71 121 72 
<< m1 >>
rect 121 71 122 72 
<< pdiffusion >>
rect 121 71 122 72 
<< pdiffusion >>
rect 122 71 123 72 
<< pdiffusion >>
rect 123 71 124 72 
<< pdiffusion >>
rect 124 71 125 72 
<< pdiffusion >>
rect 125 71 126 72 
<< m1 >>
rect 127 71 128 72 
<< m1 >>
rect 129 71 130 72 
<< pdiffusion >>
rect 138 71 139 72 
<< pdiffusion >>
rect 139 71 140 72 
<< pdiffusion >>
rect 140 71 141 72 
<< pdiffusion >>
rect 141 71 142 72 
<< m1 >>
rect 142 71 143 72 
<< pdiffusion >>
rect 142 71 143 72 
<< pdiffusion >>
rect 143 71 144 72 
<< m1 >>
rect 145 71 146 72 
<< m1 >>
rect 10 72 11 73 
<< m1 >>
rect 13 72 14 73 
<< m1 >>
rect 16 72 17 73 
<< m2 >>
rect 24 72 25 73 
<< m1 >>
rect 28 72 29 73 
<< m1 >>
rect 34 72 35 73 
<< m1 >>
rect 49 72 50 73 
<< m1 >>
rect 52 72 53 73 
<< m1 >>
rect 55 72 56 73 
<< m2 >>
rect 55 72 56 73 
<< m1 >>
rect 57 72 58 73 
<< m2 >>
rect 63 72 64 73 
<< m1 >>
rect 64 72 65 73 
<< m1 >>
rect 88 72 89 73 
<< m1 >>
rect 98 72 99 73 
<< m1 >>
rect 100 72 101 73 
<< m1 >>
rect 103 72 104 73 
<< m1 >>
rect 118 72 119 73 
<< m1 >>
rect 121 72 122 73 
<< m1 >>
rect 127 72 128 73 
<< m1 >>
rect 129 72 130 73 
<< m1 >>
rect 142 72 143 73 
<< m1 >>
rect 145 72 146 73 
<< m1 >>
rect 10 73 11 74 
<< m1 >>
rect 11 73 12 74 
<< m1 >>
rect 12 73 13 74 
<< m1 >>
rect 13 73 14 74 
<< m1 >>
rect 16 73 17 74 
<< m1 >>
rect 17 73 18 74 
<< m1 >>
rect 18 73 19 74 
<< m1 >>
rect 19 73 20 74 
<< m1 >>
rect 20 73 21 74 
<< m1 >>
rect 21 73 22 74 
<< m1 >>
rect 22 73 23 74 
<< m1 >>
rect 23 73 24 74 
<< m1 >>
rect 24 73 25 74 
<< m2 >>
rect 24 73 25 74 
<< m1 >>
rect 25 73 26 74 
<< m1 >>
rect 26 73 27 74 
<< m2 >>
rect 26 73 27 74 
<< m2c >>
rect 26 73 27 74 
<< m1 >>
rect 26 73 27 74 
<< m2 >>
rect 26 73 27 74 
<< m2 >>
rect 27 73 28 74 
<< m1 >>
rect 28 73 29 74 
<< m2 >>
rect 28 73 29 74 
<< m2 >>
rect 29 73 30 74 
<< m1 >>
rect 30 73 31 74 
<< m2 >>
rect 30 73 31 74 
<< m2c >>
rect 30 73 31 74 
<< m1 >>
rect 30 73 31 74 
<< m2 >>
rect 30 73 31 74 
<< m1 >>
rect 34 73 35 74 
<< m1 >>
rect 35 73 36 74 
<< m1 >>
rect 36 73 37 74 
<< m1 >>
rect 37 73 38 74 
<< m1 >>
rect 46 73 47 74 
<< m1 >>
rect 47 73 48 74 
<< m1 >>
rect 48 73 49 74 
<< m1 >>
rect 49 73 50 74 
<< m1 >>
rect 52 73 53 74 
<< m1 >>
rect 53 73 54 74 
<< m2 >>
rect 53 73 54 74 
<< m2c >>
rect 53 73 54 74 
<< m1 >>
rect 53 73 54 74 
<< m2 >>
rect 53 73 54 74 
<< m2 >>
rect 54 73 55 74 
<< m1 >>
rect 55 73 56 74 
<< m2 >>
rect 55 73 56 74 
<< m1 >>
rect 57 73 58 74 
<< m2 >>
rect 63 73 64 74 
<< m1 >>
rect 64 73 65 74 
<< m2 >>
rect 64 73 65 74 
<< m2 >>
rect 65 73 66 74 
<< m1 >>
rect 66 73 67 74 
<< m2 >>
rect 66 73 67 74 
<< m2c >>
rect 66 73 67 74 
<< m1 >>
rect 66 73 67 74 
<< m2 >>
rect 66 73 67 74 
<< m1 >>
rect 88 73 89 74 
<< m1 >>
rect 98 73 99 74 
<< m1 >>
rect 100 73 101 74 
<< m1 >>
rect 103 73 104 74 
<< m1 >>
rect 118 73 119 74 
<< m1 >>
rect 121 73 122 74 
<< m1 >>
rect 127 73 128 74 
<< m1 >>
rect 129 73 130 74 
<< m1 >>
rect 142 73 143 74 
<< m1 >>
rect 145 73 146 74 
<< m2 >>
rect 24 74 25 75 
<< m1 >>
rect 28 74 29 75 
<< m1 >>
rect 30 74 31 75 
<< m2 >>
rect 33 74 34 75 
<< m2 >>
rect 34 74 35 75 
<< m2 >>
rect 35 74 36 75 
<< m2 >>
rect 36 74 37 75 
<< m1 >>
rect 37 74 38 75 
<< m2 >>
rect 37 74 38 75 
<< m2 >>
rect 38 74 39 75 
<< m1 >>
rect 39 74 40 75 
<< m2 >>
rect 39 74 40 75 
<< m2c >>
rect 39 74 40 75 
<< m1 >>
rect 39 74 40 75 
<< m2 >>
rect 39 74 40 75 
<< m1 >>
rect 46 74 47 75 
<< m1 >>
rect 55 74 56 75 
<< m1 >>
rect 57 74 58 75 
<< m1 >>
rect 64 74 65 75 
<< m1 >>
rect 66 74 67 75 
<< m1 >>
rect 88 74 89 75 
<< m2 >>
rect 88 74 89 75 
<< m2c >>
rect 88 74 89 75 
<< m1 >>
rect 88 74 89 75 
<< m2 >>
rect 88 74 89 75 
<< m1 >>
rect 98 74 99 75 
<< m1 >>
rect 100 74 101 75 
<< m2 >>
rect 100 74 101 75 
<< m2c >>
rect 100 74 101 75 
<< m1 >>
rect 100 74 101 75 
<< m2 >>
rect 100 74 101 75 
<< m1 >>
rect 103 74 104 75 
<< m1 >>
rect 104 74 105 75 
<< m1 >>
rect 105 74 106 75 
<< m1 >>
rect 106 74 107 75 
<< m1 >>
rect 107 74 108 75 
<< m1 >>
rect 108 74 109 75 
<< m1 >>
rect 109 74 110 75 
<< m1 >>
rect 110 74 111 75 
<< m1 >>
rect 111 74 112 75 
<< m1 >>
rect 112 74 113 75 
<< m1 >>
rect 113 74 114 75 
<< m1 >>
rect 114 74 115 75 
<< m1 >>
rect 115 74 116 75 
<< m1 >>
rect 116 74 117 75 
<< m2 >>
rect 116 74 117 75 
<< m2c >>
rect 116 74 117 75 
<< m1 >>
rect 116 74 117 75 
<< m2 >>
rect 116 74 117 75 
<< m2 >>
rect 117 74 118 75 
<< m1 >>
rect 118 74 119 75 
<< m2 >>
rect 118 74 119 75 
<< m2 >>
rect 119 74 120 75 
<< m2 >>
rect 120 74 121 75 
<< m1 >>
rect 121 74 122 75 
<< m1 >>
rect 127 74 128 75 
<< m2 >>
rect 127 74 128 75 
<< m2c >>
rect 127 74 128 75 
<< m1 >>
rect 127 74 128 75 
<< m2 >>
rect 127 74 128 75 
<< m1 >>
rect 129 74 130 75 
<< m2 >>
rect 129 74 130 75 
<< m2c >>
rect 129 74 130 75 
<< m1 >>
rect 129 74 130 75 
<< m2 >>
rect 129 74 130 75 
<< m1 >>
rect 142 74 143 75 
<< m1 >>
rect 145 74 146 75 
<< m1 >>
rect 24 75 25 76 
<< m2 >>
rect 24 75 25 76 
<< m2c >>
rect 24 75 25 76 
<< m1 >>
rect 24 75 25 76 
<< m2 >>
rect 24 75 25 76 
<< m1 >>
rect 28 75 29 76 
<< m1 >>
rect 30 75 31 76 
<< m2 >>
rect 33 75 34 76 
<< m1 >>
rect 37 75 38 76 
<< m1 >>
rect 39 75 40 76 
<< m1 >>
rect 46 75 47 76 
<< m1 >>
rect 55 75 56 76 
<< m1 >>
rect 57 75 58 76 
<< m1 >>
rect 64 75 65 76 
<< m1 >>
rect 66 75 67 76 
<< m2 >>
rect 88 75 89 76 
<< m1 >>
rect 98 75 99 76 
<< m2 >>
rect 100 75 101 76 
<< m1 >>
rect 118 75 119 76 
<< m2 >>
rect 120 75 121 76 
<< m1 >>
rect 121 75 122 76 
<< m2 >>
rect 127 75 128 76 
<< m2 >>
rect 129 75 130 76 
<< m1 >>
rect 142 75 143 76 
<< m1 >>
rect 145 75 146 76 
<< m1 >>
rect 10 76 11 77 
<< m1 >>
rect 11 76 12 77 
<< m1 >>
rect 12 76 13 77 
<< m1 >>
rect 13 76 14 77 
<< m1 >>
rect 14 76 15 77 
<< m1 >>
rect 15 76 16 77 
<< m1 >>
rect 16 76 17 77 
<< m1 >>
rect 17 76 18 77 
<< m1 >>
rect 18 76 19 77 
<< m1 >>
rect 19 76 20 77 
<< m1 >>
rect 20 76 21 77 
<< m1 >>
rect 21 76 22 77 
<< m1 >>
rect 22 76 23 77 
<< m1 >>
rect 23 76 24 77 
<< m1 >>
rect 24 76 25 77 
<< m1 >>
rect 28 76 29 77 
<< m1 >>
rect 30 76 31 77 
<< m1 >>
rect 31 76 32 77 
<< m1 >>
rect 32 76 33 77 
<< m1 >>
rect 33 76 34 77 
<< m2 >>
rect 33 76 34 77 
<< m1 >>
rect 34 76 35 77 
<< m1 >>
rect 35 76 36 77 
<< m2 >>
rect 35 76 36 77 
<< m2c >>
rect 35 76 36 77 
<< m1 >>
rect 35 76 36 77 
<< m2 >>
rect 35 76 36 77 
<< m2 >>
rect 36 76 37 77 
<< m1 >>
rect 37 76 38 77 
<< m2 >>
rect 37 76 38 77 
<< m1 >>
rect 39 76 40 77 
<< m1 >>
rect 46 76 47 77 
<< m1 >>
rect 55 76 56 77 
<< m1 >>
rect 57 76 58 77 
<< m1 >>
rect 60 76 61 77 
<< m1 >>
rect 61 76 62 77 
<< m1 >>
rect 62 76 63 77 
<< m2 >>
rect 62 76 63 77 
<< m2c >>
rect 62 76 63 77 
<< m1 >>
rect 62 76 63 77 
<< m2 >>
rect 62 76 63 77 
<< m2 >>
rect 63 76 64 77 
<< m1 >>
rect 64 76 65 77 
<< m2 >>
rect 64 76 65 77 
<< m2 >>
rect 65 76 66 77 
<< m1 >>
rect 66 76 67 77 
<< m2 >>
rect 66 76 67 77 
<< m1 >>
rect 67 76 68 77 
<< m2 >>
rect 67 76 68 77 
<< m1 >>
rect 68 76 69 77 
<< m2 >>
rect 68 76 69 77 
<< m1 >>
rect 69 76 70 77 
<< m2 >>
rect 69 76 70 77 
<< m1 >>
rect 70 76 71 77 
<< m2 >>
rect 70 76 71 77 
<< m1 >>
rect 71 76 72 77 
<< m2 >>
rect 71 76 72 77 
<< m1 >>
rect 72 76 73 77 
<< m2 >>
rect 72 76 73 77 
<< m1 >>
rect 73 76 74 77 
<< m2 >>
rect 73 76 74 77 
<< m1 >>
rect 74 76 75 77 
<< m2 >>
rect 74 76 75 77 
<< m1 >>
rect 75 76 76 77 
<< m2 >>
rect 75 76 76 77 
<< m1 >>
rect 76 76 77 77 
<< m2 >>
rect 76 76 77 77 
<< m1 >>
rect 77 76 78 77 
<< m2 >>
rect 77 76 78 77 
<< m1 >>
rect 78 76 79 77 
<< m2 >>
rect 78 76 79 77 
<< m1 >>
rect 79 76 80 77 
<< m2 >>
rect 79 76 80 77 
<< m1 >>
rect 80 76 81 77 
<< m2 >>
rect 80 76 81 77 
<< m1 >>
rect 81 76 82 77 
<< m2 >>
rect 81 76 82 77 
<< m1 >>
rect 82 76 83 77 
<< m2 >>
rect 82 76 83 77 
<< m1 >>
rect 83 76 84 77 
<< m2 >>
rect 83 76 84 77 
<< m1 >>
rect 84 76 85 77 
<< m2 >>
rect 84 76 85 77 
<< m1 >>
rect 85 76 86 77 
<< m2 >>
rect 85 76 86 77 
<< m1 >>
rect 86 76 87 77 
<< m2 >>
rect 86 76 87 77 
<< m1 >>
rect 87 76 88 77 
<< m2 >>
rect 87 76 88 77 
<< m1 >>
rect 88 76 89 77 
<< m2 >>
rect 88 76 89 77 
<< m1 >>
rect 89 76 90 77 
<< m1 >>
rect 90 76 91 77 
<< m1 >>
rect 91 76 92 77 
<< m1 >>
rect 98 76 99 77 
<< m1 >>
rect 100 76 101 77 
<< m2 >>
rect 100 76 101 77 
<< m1 >>
rect 101 76 102 77 
<< m1 >>
rect 102 76 103 77 
<< m1 >>
rect 103 76 104 77 
<< m1 >>
rect 104 76 105 77 
<< m1 >>
rect 105 76 106 77 
<< m1 >>
rect 106 76 107 77 
<< m1 >>
rect 107 76 108 77 
<< m1 >>
rect 108 76 109 77 
<< m1 >>
rect 109 76 110 77 
<< m1 >>
rect 110 76 111 77 
<< m1 >>
rect 111 76 112 77 
<< m1 >>
rect 112 76 113 77 
<< m1 >>
rect 113 76 114 77 
<< m1 >>
rect 114 76 115 77 
<< m1 >>
rect 115 76 116 77 
<< m1 >>
rect 116 76 117 77 
<< m1 >>
rect 117 76 118 77 
<< m1 >>
rect 118 76 119 77 
<< m2 >>
rect 120 76 121 77 
<< m1 >>
rect 121 76 122 77 
<< m1 >>
rect 122 76 123 77 
<< m1 >>
rect 123 76 124 77 
<< m1 >>
rect 124 76 125 77 
<< m1 >>
rect 125 76 126 77 
<< m1 >>
rect 126 76 127 77 
<< m1 >>
rect 127 76 128 77 
<< m2 >>
rect 127 76 128 77 
<< m1 >>
rect 128 76 129 77 
<< m1 >>
rect 129 76 130 77 
<< m2 >>
rect 129 76 130 77 
<< m1 >>
rect 130 76 131 77 
<< m1 >>
rect 131 76 132 77 
<< m1 >>
rect 132 76 133 77 
<< m1 >>
rect 133 76 134 77 
<< m1 >>
rect 134 76 135 77 
<< m1 >>
rect 135 76 136 77 
<< m1 >>
rect 136 76 137 77 
<< m1 >>
rect 137 76 138 77 
<< m1 >>
rect 138 76 139 77 
<< m1 >>
rect 139 76 140 77 
<< m1 >>
rect 140 76 141 77 
<< m1 >>
rect 141 76 142 77 
<< m1 >>
rect 142 76 143 77 
<< m1 >>
rect 145 76 146 77 
<< m1 >>
rect 10 77 11 78 
<< m1 >>
rect 28 77 29 78 
<< m2 >>
rect 33 77 34 78 
<< m1 >>
rect 37 77 38 78 
<< m2 >>
rect 37 77 38 78 
<< m1 >>
rect 39 77 40 78 
<< m1 >>
rect 46 77 47 78 
<< m1 >>
rect 55 77 56 78 
<< m1 >>
rect 57 77 58 78 
<< m1 >>
rect 60 77 61 78 
<< m1 >>
rect 64 77 65 78 
<< m1 >>
rect 91 77 92 78 
<< m1 >>
rect 98 77 99 78 
<< m1 >>
rect 100 77 101 78 
<< m2 >>
rect 100 77 101 78 
<< m2 >>
rect 120 77 121 78 
<< m2 >>
rect 121 77 122 78 
<< m2 >>
rect 122 77 123 78 
<< m2 >>
rect 123 77 124 78 
<< m2 >>
rect 124 77 125 78 
<< m2 >>
rect 125 77 126 78 
<< m2 >>
rect 127 77 128 78 
<< m2 >>
rect 129 77 130 78 
<< m1 >>
rect 145 77 146 78 
<< m1 >>
rect 10 78 11 79 
<< m1 >>
rect 28 78 29 79 
<< m1 >>
rect 33 78 34 79 
<< m2 >>
rect 33 78 34 79 
<< m2c >>
rect 33 78 34 79 
<< m1 >>
rect 33 78 34 79 
<< m2 >>
rect 33 78 34 79 
<< m1 >>
rect 34 78 35 79 
<< m1 >>
rect 37 78 38 79 
<< m2 >>
rect 37 78 38 79 
<< m1 >>
rect 39 78 40 79 
<< m2 >>
rect 39 78 40 79 
<< m2c >>
rect 39 78 40 79 
<< m1 >>
rect 39 78 40 79 
<< m2 >>
rect 39 78 40 79 
<< m1 >>
rect 46 78 47 79 
<< m1 >>
rect 55 78 56 79 
<< m1 >>
rect 57 78 58 79 
<< m1 >>
rect 60 78 61 79 
<< m1 >>
rect 64 78 65 79 
<< m1 >>
rect 91 78 92 79 
<< m1 >>
rect 98 78 99 79 
<< m1 >>
rect 100 78 101 79 
<< m2 >>
rect 100 78 101 79 
<< m2 >>
rect 101 78 102 79 
<< m1 >>
rect 102 78 103 79 
<< m2 >>
rect 102 78 103 79 
<< m2c >>
rect 102 78 103 79 
<< m1 >>
rect 102 78 103 79 
<< m2 >>
rect 102 78 103 79 
<< m1 >>
rect 103 78 104 79 
<< m1 >>
rect 125 78 126 79 
<< m2 >>
rect 125 78 126 79 
<< m2c >>
rect 125 78 126 79 
<< m1 >>
rect 125 78 126 79 
<< m2 >>
rect 125 78 126 79 
<< m1 >>
rect 127 78 128 79 
<< m2 >>
rect 127 78 128 79 
<< m2c >>
rect 127 78 128 79 
<< m1 >>
rect 127 78 128 79 
<< m2 >>
rect 127 78 128 79 
<< m1 >>
rect 129 78 130 79 
<< m2 >>
rect 129 78 130 79 
<< m2c >>
rect 129 78 130 79 
<< m1 >>
rect 129 78 130 79 
<< m2 >>
rect 129 78 130 79 
<< m1 >>
rect 145 78 146 79 
<< m1 >>
rect 10 79 11 80 
<< m1 >>
rect 28 79 29 80 
<< m1 >>
rect 34 79 35 80 
<< m1 >>
rect 37 79 38 80 
<< m2 >>
rect 37 79 38 80 
<< m2 >>
rect 39 79 40 80 
<< m2 >>
rect 45 79 46 80 
<< m1 >>
rect 46 79 47 80 
<< m2 >>
rect 46 79 47 80 
<< m2 >>
rect 47 79 48 80 
<< m1 >>
rect 48 79 49 80 
<< m2 >>
rect 48 79 49 80 
<< m1 >>
rect 49 79 50 80 
<< m2 >>
rect 49 79 50 80 
<< m1 >>
rect 50 79 51 80 
<< m2 >>
rect 50 79 51 80 
<< m1 >>
rect 51 79 52 80 
<< m1 >>
rect 52 79 53 80 
<< m1 >>
rect 53 79 54 80 
<< m2 >>
rect 53 79 54 80 
<< m2c >>
rect 53 79 54 80 
<< m1 >>
rect 53 79 54 80 
<< m2 >>
rect 53 79 54 80 
<< m2 >>
rect 54 79 55 80 
<< m1 >>
rect 55 79 56 80 
<< m2 >>
rect 55 79 56 80 
<< m2 >>
rect 56 79 57 80 
<< m1 >>
rect 57 79 58 80 
<< m2 >>
rect 57 79 58 80 
<< m2c >>
rect 57 79 58 80 
<< m1 >>
rect 57 79 58 80 
<< m2 >>
rect 57 79 58 80 
<< m1 >>
rect 60 79 61 80 
<< m2 >>
rect 63 79 64 80 
<< m1 >>
rect 64 79 65 80 
<< m2 >>
rect 64 79 65 80 
<< m2 >>
rect 65 79 66 80 
<< m1 >>
rect 66 79 67 80 
<< m2 >>
rect 66 79 67 80 
<< m2c >>
rect 66 79 67 80 
<< m1 >>
rect 66 79 67 80 
<< m2 >>
rect 66 79 67 80 
<< m1 >>
rect 67 79 68 80 
<< m1 >>
rect 68 79 69 80 
<< m2 >>
rect 68 79 69 80 
<< m2c >>
rect 68 79 69 80 
<< m1 >>
rect 68 79 69 80 
<< m2 >>
rect 68 79 69 80 
<< m1 >>
rect 91 79 92 80 
<< m1 >>
rect 98 79 99 80 
<< m1 >>
rect 100 79 101 80 
<< m1 >>
rect 103 79 104 80 
<< m1 >>
rect 125 79 126 80 
<< m1 >>
rect 127 79 128 80 
<< m1 >>
rect 129 79 130 80 
<< m1 >>
rect 145 79 146 80 
<< m1 >>
rect 10 80 11 81 
<< m1 >>
rect 28 80 29 81 
<< m1 >>
rect 34 80 35 81 
<< m1 >>
rect 37 80 38 81 
<< m2 >>
rect 37 80 38 81 
<< m2 >>
rect 39 80 40 81 
<< m1 >>
rect 40 80 41 81 
<< m1 >>
rect 41 80 42 81 
<< m1 >>
rect 42 80 43 81 
<< m1 >>
rect 43 80 44 81 
<< m1 >>
rect 44 80 45 81 
<< m2 >>
rect 44 80 45 81 
<< m2c >>
rect 44 80 45 81 
<< m1 >>
rect 44 80 45 81 
<< m2 >>
rect 44 80 45 81 
<< m2 >>
rect 45 80 46 81 
<< m1 >>
rect 46 80 47 81 
<< m1 >>
rect 48 80 49 81 
<< m2 >>
rect 50 80 51 81 
<< m1 >>
rect 55 80 56 81 
<< m1 >>
rect 60 80 61 81 
<< m2 >>
rect 63 80 64 81 
<< m1 >>
rect 64 80 65 81 
<< m2 >>
rect 68 80 69 81 
<< m2 >>
rect 69 80 70 81 
<< m2 >>
rect 70 80 71 81 
<< m1 >>
rect 91 80 92 81 
<< m1 >>
rect 98 80 99 81 
<< m1 >>
rect 100 80 101 81 
<< m1 >>
rect 103 80 104 81 
<< m1 >>
rect 125 80 126 81 
<< m2 >>
rect 125 80 126 81 
<< m2c >>
rect 125 80 126 81 
<< m1 >>
rect 125 80 126 81 
<< m2 >>
rect 125 80 126 81 
<< m2 >>
rect 126 80 127 81 
<< m1 >>
rect 127 80 128 81 
<< m2 >>
rect 127 80 128 81 
<< m2 >>
rect 128 80 129 81 
<< m1 >>
rect 129 80 130 81 
<< m2 >>
rect 129 80 130 81 
<< m2c >>
rect 129 80 130 81 
<< m1 >>
rect 129 80 130 81 
<< m2 >>
rect 129 80 130 81 
<< m1 >>
rect 145 80 146 81 
<< m1 >>
rect 10 81 11 82 
<< m1 >>
rect 28 81 29 82 
<< m1 >>
rect 34 81 35 82 
<< m1 >>
rect 37 81 38 82 
<< m2 >>
rect 37 81 38 82 
<< m2 >>
rect 39 81 40 82 
<< m1 >>
rect 40 81 41 82 
<< m1 >>
rect 46 81 47 82 
<< m1 >>
rect 48 81 49 82 
<< m1 >>
rect 50 81 51 82 
<< m2 >>
rect 50 81 51 82 
<< m2c >>
rect 50 81 51 82 
<< m1 >>
rect 50 81 51 82 
<< m2 >>
rect 50 81 51 82 
<< m1 >>
rect 51 81 52 82 
<< m1 >>
rect 52 81 53 82 
<< m1 >>
rect 55 81 56 82 
<< m1 >>
rect 60 81 61 82 
<< m2 >>
rect 63 81 64 82 
<< m1 >>
rect 64 81 65 82 
<< m1 >>
rect 67 81 68 82 
<< m1 >>
rect 68 81 69 82 
<< m1 >>
rect 69 81 70 82 
<< m1 >>
rect 70 81 71 82 
<< m2 >>
rect 70 81 71 82 
<< m1 >>
rect 71 81 72 82 
<< m1 >>
rect 72 81 73 82 
<< m1 >>
rect 73 81 74 82 
<< m1 >>
rect 74 81 75 82 
<< m1 >>
rect 75 81 76 82 
<< m1 >>
rect 76 81 77 82 
<< m1 >>
rect 77 81 78 82 
<< m1 >>
rect 78 81 79 82 
<< m1 >>
rect 79 81 80 82 
<< m1 >>
rect 80 81 81 82 
<< m1 >>
rect 81 81 82 82 
<< m1 >>
rect 82 81 83 82 
<< m1 >>
rect 91 81 92 82 
<< m1 >>
rect 98 81 99 82 
<< m1 >>
rect 100 81 101 82 
<< m1 >>
rect 103 81 104 82 
<< m1 >>
rect 127 81 128 82 
<< m1 >>
rect 145 81 146 82 
<< m1 >>
rect 10 82 11 83 
<< m2 >>
rect 27 82 28 83 
<< m1 >>
rect 28 82 29 83 
<< m2 >>
rect 28 82 29 83 
<< m2 >>
rect 29 82 30 83 
<< m1 >>
rect 30 82 31 83 
<< m2 >>
rect 30 82 31 83 
<< m2c >>
rect 30 82 31 83 
<< m1 >>
rect 30 82 31 83 
<< m2 >>
rect 30 82 31 83 
<< m1 >>
rect 31 82 32 83 
<< m1 >>
rect 34 82 35 83 
<< m1 >>
rect 37 82 38 83 
<< m2 >>
rect 37 82 38 83 
<< m2 >>
rect 39 82 40 83 
<< m1 >>
rect 40 82 41 83 
<< m2 >>
rect 45 82 46 83 
<< m1 >>
rect 46 82 47 83 
<< m2 >>
rect 46 82 47 83 
<< m2 >>
rect 47 82 48 83 
<< m1 >>
rect 48 82 49 83 
<< m2 >>
rect 48 82 49 83 
<< m2c >>
rect 48 82 49 83 
<< m1 >>
rect 48 82 49 83 
<< m2 >>
rect 48 82 49 83 
<< m1 >>
rect 52 82 53 83 
<< m1 >>
rect 55 82 56 83 
<< m1 >>
rect 60 82 61 83 
<< m2 >>
rect 63 82 64 83 
<< m1 >>
rect 64 82 65 83 
<< m1 >>
rect 67 82 68 83 
<< m2 >>
rect 70 82 71 83 
<< m1 >>
rect 82 82 83 83 
<< m1 >>
rect 91 82 92 83 
<< m1 >>
rect 98 82 99 83 
<< m1 >>
rect 100 82 101 83 
<< m1 >>
rect 103 82 104 83 
<< m1 >>
rect 106 82 107 83 
<< m1 >>
rect 107 82 108 83 
<< m1 >>
rect 108 82 109 83 
<< m1 >>
rect 109 82 110 83 
<< m1 >>
rect 127 82 128 83 
<< m1 >>
rect 145 82 146 83 
<< m1 >>
rect 10 83 11 84 
<< m2 >>
rect 27 83 28 84 
<< m1 >>
rect 28 83 29 84 
<< m1 >>
rect 31 83 32 84 
<< m1 >>
rect 34 83 35 84 
<< m1 >>
rect 37 83 38 84 
<< m2 >>
rect 37 83 38 84 
<< m2 >>
rect 39 83 40 84 
<< m1 >>
rect 40 83 41 84 
<< m2 >>
rect 45 83 46 84 
<< m1 >>
rect 46 83 47 84 
<< m1 >>
rect 52 83 53 84 
<< m1 >>
rect 55 83 56 84 
<< m1 >>
rect 60 83 61 84 
<< m2 >>
rect 63 83 64 84 
<< m1 >>
rect 64 83 65 84 
<< m1 >>
rect 67 83 68 84 
<< m1 >>
rect 70 83 71 84 
<< m2 >>
rect 70 83 71 84 
<< m2c >>
rect 70 83 71 84 
<< m1 >>
rect 70 83 71 84 
<< m2 >>
rect 70 83 71 84 
<< m1 >>
rect 82 83 83 84 
<< m1 >>
rect 91 83 92 84 
<< m1 >>
rect 98 83 99 84 
<< m1 >>
rect 100 83 101 84 
<< m1 >>
rect 103 83 104 84 
<< m1 >>
rect 106 83 107 84 
<< m1 >>
rect 109 83 110 84 
<< m1 >>
rect 127 83 128 84 
<< m1 >>
rect 145 83 146 84 
<< m1 >>
rect 10 84 11 85 
<< pdiffusion >>
rect 12 84 13 85 
<< pdiffusion >>
rect 13 84 14 85 
<< pdiffusion >>
rect 14 84 15 85 
<< pdiffusion >>
rect 15 84 16 85 
<< pdiffusion >>
rect 16 84 17 85 
<< pdiffusion >>
rect 17 84 18 85 
<< m2 >>
rect 27 84 28 85 
<< m1 >>
rect 28 84 29 85 
<< pdiffusion >>
rect 30 84 31 85 
<< m1 >>
rect 31 84 32 85 
<< pdiffusion >>
rect 31 84 32 85 
<< pdiffusion >>
rect 32 84 33 85 
<< pdiffusion >>
rect 33 84 34 85 
<< m1 >>
rect 34 84 35 85 
<< pdiffusion >>
rect 34 84 35 85 
<< pdiffusion >>
rect 35 84 36 85 
<< m1 >>
rect 37 84 38 85 
<< m2 >>
rect 37 84 38 85 
<< m2 >>
rect 39 84 40 85 
<< m1 >>
rect 40 84 41 85 
<< m2 >>
rect 45 84 46 85 
<< m1 >>
rect 46 84 47 85 
<< pdiffusion >>
rect 48 84 49 85 
<< pdiffusion >>
rect 49 84 50 85 
<< pdiffusion >>
rect 50 84 51 85 
<< pdiffusion >>
rect 51 84 52 85 
<< m1 >>
rect 52 84 53 85 
<< pdiffusion >>
rect 52 84 53 85 
<< pdiffusion >>
rect 53 84 54 85 
<< m1 >>
rect 55 84 56 85 
<< m1 >>
rect 60 84 61 85 
<< m2 >>
rect 63 84 64 85 
<< m1 >>
rect 64 84 65 85 
<< pdiffusion >>
rect 66 84 67 85 
<< m1 >>
rect 67 84 68 85 
<< pdiffusion >>
rect 67 84 68 85 
<< pdiffusion >>
rect 68 84 69 85 
<< pdiffusion >>
rect 69 84 70 85 
<< m1 >>
rect 70 84 71 85 
<< pdiffusion >>
rect 70 84 71 85 
<< pdiffusion >>
rect 71 84 72 85 
<< m1 >>
rect 82 84 83 85 
<< pdiffusion >>
rect 84 84 85 85 
<< pdiffusion >>
rect 85 84 86 85 
<< pdiffusion >>
rect 86 84 87 85 
<< pdiffusion >>
rect 87 84 88 85 
<< pdiffusion >>
rect 88 84 89 85 
<< pdiffusion >>
rect 89 84 90 85 
<< m1 >>
rect 91 84 92 85 
<< m1 >>
rect 98 84 99 85 
<< m1 >>
rect 100 84 101 85 
<< pdiffusion >>
rect 102 84 103 85 
<< m1 >>
rect 103 84 104 85 
<< pdiffusion >>
rect 103 84 104 85 
<< pdiffusion >>
rect 104 84 105 85 
<< pdiffusion >>
rect 105 84 106 85 
<< m1 >>
rect 106 84 107 85 
<< pdiffusion >>
rect 106 84 107 85 
<< pdiffusion >>
rect 107 84 108 85 
<< m1 >>
rect 109 84 110 85 
<< m1 >>
rect 127 84 128 85 
<< pdiffusion >>
rect 138 84 139 85 
<< pdiffusion >>
rect 139 84 140 85 
<< pdiffusion >>
rect 140 84 141 85 
<< pdiffusion >>
rect 141 84 142 85 
<< pdiffusion >>
rect 142 84 143 85 
<< pdiffusion >>
rect 143 84 144 85 
<< m1 >>
rect 145 84 146 85 
<< m1 >>
rect 10 85 11 86 
<< pdiffusion >>
rect 12 85 13 86 
<< pdiffusion >>
rect 13 85 14 86 
<< pdiffusion >>
rect 14 85 15 86 
<< pdiffusion >>
rect 15 85 16 86 
<< pdiffusion >>
rect 16 85 17 86 
<< pdiffusion >>
rect 17 85 18 86 
<< m2 >>
rect 27 85 28 86 
<< m1 >>
rect 28 85 29 86 
<< pdiffusion >>
rect 30 85 31 86 
<< pdiffusion >>
rect 31 85 32 86 
<< pdiffusion >>
rect 32 85 33 86 
<< pdiffusion >>
rect 33 85 34 86 
<< pdiffusion >>
rect 34 85 35 86 
<< pdiffusion >>
rect 35 85 36 86 
<< m1 >>
rect 37 85 38 86 
<< m2 >>
rect 37 85 38 86 
<< m2 >>
rect 39 85 40 86 
<< m1 >>
rect 40 85 41 86 
<< m2 >>
rect 45 85 46 86 
<< m1 >>
rect 46 85 47 86 
<< pdiffusion >>
rect 48 85 49 86 
<< pdiffusion >>
rect 49 85 50 86 
<< pdiffusion >>
rect 50 85 51 86 
<< pdiffusion >>
rect 51 85 52 86 
<< pdiffusion >>
rect 52 85 53 86 
<< pdiffusion >>
rect 53 85 54 86 
<< m1 >>
rect 55 85 56 86 
<< m1 >>
rect 60 85 61 86 
<< m2 >>
rect 63 85 64 86 
<< m1 >>
rect 64 85 65 86 
<< pdiffusion >>
rect 66 85 67 86 
<< pdiffusion >>
rect 67 85 68 86 
<< pdiffusion >>
rect 68 85 69 86 
<< pdiffusion >>
rect 69 85 70 86 
<< pdiffusion >>
rect 70 85 71 86 
<< pdiffusion >>
rect 71 85 72 86 
<< m1 >>
rect 82 85 83 86 
<< pdiffusion >>
rect 84 85 85 86 
<< pdiffusion >>
rect 85 85 86 86 
<< pdiffusion >>
rect 86 85 87 86 
<< pdiffusion >>
rect 87 85 88 86 
<< pdiffusion >>
rect 88 85 89 86 
<< pdiffusion >>
rect 89 85 90 86 
<< m1 >>
rect 91 85 92 86 
<< m1 >>
rect 98 85 99 86 
<< m1 >>
rect 100 85 101 86 
<< pdiffusion >>
rect 102 85 103 86 
<< pdiffusion >>
rect 103 85 104 86 
<< pdiffusion >>
rect 104 85 105 86 
<< pdiffusion >>
rect 105 85 106 86 
<< pdiffusion >>
rect 106 85 107 86 
<< pdiffusion >>
rect 107 85 108 86 
<< m1 >>
rect 109 85 110 86 
<< m1 >>
rect 127 85 128 86 
<< pdiffusion >>
rect 138 85 139 86 
<< pdiffusion >>
rect 139 85 140 86 
<< pdiffusion >>
rect 140 85 141 86 
<< pdiffusion >>
rect 141 85 142 86 
<< pdiffusion >>
rect 142 85 143 86 
<< pdiffusion >>
rect 143 85 144 86 
<< m1 >>
rect 145 85 146 86 
<< m1 >>
rect 10 86 11 87 
<< pdiffusion >>
rect 12 86 13 87 
<< pdiffusion >>
rect 13 86 14 87 
<< pdiffusion >>
rect 14 86 15 87 
<< pdiffusion >>
rect 15 86 16 87 
<< pdiffusion >>
rect 16 86 17 87 
<< pdiffusion >>
rect 17 86 18 87 
<< m2 >>
rect 27 86 28 87 
<< m1 >>
rect 28 86 29 87 
<< pdiffusion >>
rect 30 86 31 87 
<< pdiffusion >>
rect 31 86 32 87 
<< pdiffusion >>
rect 32 86 33 87 
<< pdiffusion >>
rect 33 86 34 87 
<< pdiffusion >>
rect 34 86 35 87 
<< pdiffusion >>
rect 35 86 36 87 
<< m1 >>
rect 37 86 38 87 
<< m2 >>
rect 37 86 38 87 
<< m2 >>
rect 39 86 40 87 
<< m1 >>
rect 40 86 41 87 
<< m2 >>
rect 45 86 46 87 
<< m1 >>
rect 46 86 47 87 
<< pdiffusion >>
rect 48 86 49 87 
<< pdiffusion >>
rect 49 86 50 87 
<< pdiffusion >>
rect 50 86 51 87 
<< pdiffusion >>
rect 51 86 52 87 
<< pdiffusion >>
rect 52 86 53 87 
<< pdiffusion >>
rect 53 86 54 87 
<< m1 >>
rect 55 86 56 87 
<< m1 >>
rect 60 86 61 87 
<< m2 >>
rect 63 86 64 87 
<< m1 >>
rect 64 86 65 87 
<< pdiffusion >>
rect 66 86 67 87 
<< pdiffusion >>
rect 67 86 68 87 
<< pdiffusion >>
rect 68 86 69 87 
<< pdiffusion >>
rect 69 86 70 87 
<< pdiffusion >>
rect 70 86 71 87 
<< pdiffusion >>
rect 71 86 72 87 
<< m1 >>
rect 82 86 83 87 
<< pdiffusion >>
rect 84 86 85 87 
<< pdiffusion >>
rect 85 86 86 87 
<< pdiffusion >>
rect 86 86 87 87 
<< pdiffusion >>
rect 87 86 88 87 
<< pdiffusion >>
rect 88 86 89 87 
<< pdiffusion >>
rect 89 86 90 87 
<< m1 >>
rect 91 86 92 87 
<< m1 >>
rect 98 86 99 87 
<< m1 >>
rect 100 86 101 87 
<< pdiffusion >>
rect 102 86 103 87 
<< pdiffusion >>
rect 103 86 104 87 
<< pdiffusion >>
rect 104 86 105 87 
<< pdiffusion >>
rect 105 86 106 87 
<< pdiffusion >>
rect 106 86 107 87 
<< pdiffusion >>
rect 107 86 108 87 
<< m1 >>
rect 109 86 110 87 
<< m1 >>
rect 127 86 128 87 
<< pdiffusion >>
rect 138 86 139 87 
<< pdiffusion >>
rect 139 86 140 87 
<< pdiffusion >>
rect 140 86 141 87 
<< pdiffusion >>
rect 141 86 142 87 
<< pdiffusion >>
rect 142 86 143 87 
<< pdiffusion >>
rect 143 86 144 87 
<< m1 >>
rect 145 86 146 87 
<< m1 >>
rect 10 87 11 88 
<< pdiffusion >>
rect 12 87 13 88 
<< pdiffusion >>
rect 13 87 14 88 
<< pdiffusion >>
rect 14 87 15 88 
<< pdiffusion >>
rect 15 87 16 88 
<< pdiffusion >>
rect 16 87 17 88 
<< pdiffusion >>
rect 17 87 18 88 
<< m2 >>
rect 27 87 28 88 
<< m1 >>
rect 28 87 29 88 
<< pdiffusion >>
rect 30 87 31 88 
<< pdiffusion >>
rect 31 87 32 88 
<< pdiffusion >>
rect 32 87 33 88 
<< pdiffusion >>
rect 33 87 34 88 
<< pdiffusion >>
rect 34 87 35 88 
<< pdiffusion >>
rect 35 87 36 88 
<< m1 >>
rect 37 87 38 88 
<< m2 >>
rect 37 87 38 88 
<< m2 >>
rect 39 87 40 88 
<< m1 >>
rect 40 87 41 88 
<< m2 >>
rect 45 87 46 88 
<< m1 >>
rect 46 87 47 88 
<< pdiffusion >>
rect 48 87 49 88 
<< pdiffusion >>
rect 49 87 50 88 
<< pdiffusion >>
rect 50 87 51 88 
<< pdiffusion >>
rect 51 87 52 88 
<< pdiffusion >>
rect 52 87 53 88 
<< pdiffusion >>
rect 53 87 54 88 
<< m1 >>
rect 55 87 56 88 
<< m1 >>
rect 60 87 61 88 
<< m2 >>
rect 63 87 64 88 
<< m1 >>
rect 64 87 65 88 
<< pdiffusion >>
rect 66 87 67 88 
<< pdiffusion >>
rect 67 87 68 88 
<< pdiffusion >>
rect 68 87 69 88 
<< pdiffusion >>
rect 69 87 70 88 
<< pdiffusion >>
rect 70 87 71 88 
<< pdiffusion >>
rect 71 87 72 88 
<< m1 >>
rect 82 87 83 88 
<< pdiffusion >>
rect 84 87 85 88 
<< pdiffusion >>
rect 85 87 86 88 
<< pdiffusion >>
rect 86 87 87 88 
<< pdiffusion >>
rect 87 87 88 88 
<< pdiffusion >>
rect 88 87 89 88 
<< pdiffusion >>
rect 89 87 90 88 
<< m1 >>
rect 91 87 92 88 
<< m1 >>
rect 98 87 99 88 
<< m1 >>
rect 100 87 101 88 
<< pdiffusion >>
rect 102 87 103 88 
<< pdiffusion >>
rect 103 87 104 88 
<< pdiffusion >>
rect 104 87 105 88 
<< pdiffusion >>
rect 105 87 106 88 
<< pdiffusion >>
rect 106 87 107 88 
<< pdiffusion >>
rect 107 87 108 88 
<< m1 >>
rect 109 87 110 88 
<< m1 >>
rect 127 87 128 88 
<< pdiffusion >>
rect 138 87 139 88 
<< pdiffusion >>
rect 139 87 140 88 
<< pdiffusion >>
rect 140 87 141 88 
<< pdiffusion >>
rect 141 87 142 88 
<< pdiffusion >>
rect 142 87 143 88 
<< pdiffusion >>
rect 143 87 144 88 
<< m1 >>
rect 145 87 146 88 
<< m1 >>
rect 10 88 11 89 
<< pdiffusion >>
rect 12 88 13 89 
<< pdiffusion >>
rect 13 88 14 89 
<< pdiffusion >>
rect 14 88 15 89 
<< pdiffusion >>
rect 15 88 16 89 
<< pdiffusion >>
rect 16 88 17 89 
<< pdiffusion >>
rect 17 88 18 89 
<< m2 >>
rect 27 88 28 89 
<< m1 >>
rect 28 88 29 89 
<< pdiffusion >>
rect 30 88 31 89 
<< pdiffusion >>
rect 31 88 32 89 
<< pdiffusion >>
rect 32 88 33 89 
<< pdiffusion >>
rect 33 88 34 89 
<< pdiffusion >>
rect 34 88 35 89 
<< pdiffusion >>
rect 35 88 36 89 
<< m1 >>
rect 37 88 38 89 
<< m2 >>
rect 37 88 38 89 
<< m2 >>
rect 39 88 40 89 
<< m1 >>
rect 40 88 41 89 
<< m2 >>
rect 45 88 46 89 
<< m1 >>
rect 46 88 47 89 
<< pdiffusion >>
rect 48 88 49 89 
<< pdiffusion >>
rect 49 88 50 89 
<< pdiffusion >>
rect 50 88 51 89 
<< pdiffusion >>
rect 51 88 52 89 
<< pdiffusion >>
rect 52 88 53 89 
<< pdiffusion >>
rect 53 88 54 89 
<< m1 >>
rect 55 88 56 89 
<< m1 >>
rect 60 88 61 89 
<< m2 >>
rect 63 88 64 89 
<< m1 >>
rect 64 88 65 89 
<< pdiffusion >>
rect 66 88 67 89 
<< pdiffusion >>
rect 67 88 68 89 
<< pdiffusion >>
rect 68 88 69 89 
<< pdiffusion >>
rect 69 88 70 89 
<< pdiffusion >>
rect 70 88 71 89 
<< pdiffusion >>
rect 71 88 72 89 
<< m1 >>
rect 82 88 83 89 
<< pdiffusion >>
rect 84 88 85 89 
<< pdiffusion >>
rect 85 88 86 89 
<< pdiffusion >>
rect 86 88 87 89 
<< pdiffusion >>
rect 87 88 88 89 
<< pdiffusion >>
rect 88 88 89 89 
<< pdiffusion >>
rect 89 88 90 89 
<< m1 >>
rect 91 88 92 89 
<< m1 >>
rect 98 88 99 89 
<< m1 >>
rect 100 88 101 89 
<< pdiffusion >>
rect 102 88 103 89 
<< pdiffusion >>
rect 103 88 104 89 
<< pdiffusion >>
rect 104 88 105 89 
<< pdiffusion >>
rect 105 88 106 89 
<< pdiffusion >>
rect 106 88 107 89 
<< pdiffusion >>
rect 107 88 108 89 
<< m1 >>
rect 109 88 110 89 
<< m1 >>
rect 127 88 128 89 
<< pdiffusion >>
rect 138 88 139 89 
<< pdiffusion >>
rect 139 88 140 89 
<< pdiffusion >>
rect 140 88 141 89 
<< pdiffusion >>
rect 141 88 142 89 
<< pdiffusion >>
rect 142 88 143 89 
<< pdiffusion >>
rect 143 88 144 89 
<< m1 >>
rect 145 88 146 89 
<< m1 >>
rect 10 89 11 90 
<< pdiffusion >>
rect 12 89 13 90 
<< m1 >>
rect 13 89 14 90 
<< pdiffusion >>
rect 13 89 14 90 
<< pdiffusion >>
rect 14 89 15 90 
<< pdiffusion >>
rect 15 89 16 90 
<< m1 >>
rect 16 89 17 90 
<< pdiffusion >>
rect 16 89 17 90 
<< pdiffusion >>
rect 17 89 18 90 
<< m2 >>
rect 27 89 28 90 
<< m1 >>
rect 28 89 29 90 
<< pdiffusion >>
rect 30 89 31 90 
<< pdiffusion >>
rect 31 89 32 90 
<< pdiffusion >>
rect 32 89 33 90 
<< pdiffusion >>
rect 33 89 34 90 
<< m1 >>
rect 34 89 35 90 
<< pdiffusion >>
rect 34 89 35 90 
<< pdiffusion >>
rect 35 89 36 90 
<< m1 >>
rect 37 89 38 90 
<< m2 >>
rect 37 89 38 90 
<< m2 >>
rect 39 89 40 90 
<< m1 >>
rect 40 89 41 90 
<< m2 >>
rect 45 89 46 90 
<< m1 >>
rect 46 89 47 90 
<< pdiffusion >>
rect 48 89 49 90 
<< m1 >>
rect 49 89 50 90 
<< pdiffusion >>
rect 49 89 50 90 
<< pdiffusion >>
rect 50 89 51 90 
<< pdiffusion >>
rect 51 89 52 90 
<< m1 >>
rect 52 89 53 90 
<< pdiffusion >>
rect 52 89 53 90 
<< pdiffusion >>
rect 53 89 54 90 
<< m1 >>
rect 55 89 56 90 
<< m1 >>
rect 60 89 61 90 
<< m2 >>
rect 63 89 64 90 
<< m1 >>
rect 64 89 65 90 
<< pdiffusion >>
rect 66 89 67 90 
<< m1 >>
rect 67 89 68 90 
<< pdiffusion >>
rect 67 89 68 90 
<< pdiffusion >>
rect 68 89 69 90 
<< pdiffusion >>
rect 69 89 70 90 
<< m1 >>
rect 70 89 71 90 
<< pdiffusion >>
rect 70 89 71 90 
<< pdiffusion >>
rect 71 89 72 90 
<< m1 >>
rect 82 89 83 90 
<< pdiffusion >>
rect 84 89 85 90 
<< m1 >>
rect 85 89 86 90 
<< pdiffusion >>
rect 85 89 86 90 
<< pdiffusion >>
rect 86 89 87 90 
<< pdiffusion >>
rect 87 89 88 90 
<< m1 >>
rect 88 89 89 90 
<< pdiffusion >>
rect 88 89 89 90 
<< pdiffusion >>
rect 89 89 90 90 
<< m1 >>
rect 91 89 92 90 
<< m2 >>
rect 91 89 92 90 
<< m2c >>
rect 91 89 92 90 
<< m1 >>
rect 91 89 92 90 
<< m2 >>
rect 91 89 92 90 
<< m1 >>
rect 98 89 99 90 
<< m2 >>
rect 98 89 99 90 
<< m2c >>
rect 98 89 99 90 
<< m1 >>
rect 98 89 99 90 
<< m2 >>
rect 98 89 99 90 
<< m2 >>
rect 99 89 100 90 
<< m1 >>
rect 100 89 101 90 
<< m2 >>
rect 100 89 101 90 
<< pdiffusion >>
rect 102 89 103 90 
<< pdiffusion >>
rect 103 89 104 90 
<< pdiffusion >>
rect 104 89 105 90 
<< pdiffusion >>
rect 105 89 106 90 
<< pdiffusion >>
rect 106 89 107 90 
<< pdiffusion >>
rect 107 89 108 90 
<< m1 >>
rect 109 89 110 90 
<< m1 >>
rect 127 89 128 90 
<< pdiffusion >>
rect 138 89 139 90 
<< m1 >>
rect 139 89 140 90 
<< pdiffusion >>
rect 139 89 140 90 
<< pdiffusion >>
rect 140 89 141 90 
<< pdiffusion >>
rect 141 89 142 90 
<< m1 >>
rect 142 89 143 90 
<< pdiffusion >>
rect 142 89 143 90 
<< pdiffusion >>
rect 143 89 144 90 
<< m1 >>
rect 145 89 146 90 
<< m1 >>
rect 10 90 11 91 
<< m1 >>
rect 13 90 14 91 
<< m1 >>
rect 16 90 17 91 
<< m2 >>
rect 27 90 28 91 
<< m1 >>
rect 28 90 29 91 
<< m1 >>
rect 34 90 35 91 
<< m1 >>
rect 37 90 38 91 
<< m2 >>
rect 37 90 38 91 
<< m2 >>
rect 39 90 40 91 
<< m1 >>
rect 40 90 41 91 
<< m2 >>
rect 45 90 46 91 
<< m1 >>
rect 46 90 47 91 
<< m1 >>
rect 49 90 50 91 
<< m1 >>
rect 52 90 53 91 
<< m1 >>
rect 55 90 56 91 
<< m1 >>
rect 60 90 61 91 
<< m2 >>
rect 63 90 64 91 
<< m1 >>
rect 64 90 65 91 
<< m1 >>
rect 67 90 68 91 
<< m1 >>
rect 70 90 71 91 
<< m2 >>
rect 70 90 71 91 
<< m2c >>
rect 70 90 71 91 
<< m1 >>
rect 70 90 71 91 
<< m2 >>
rect 70 90 71 91 
<< m1 >>
rect 82 90 83 91 
<< m2 >>
rect 82 90 83 91 
<< m2c >>
rect 82 90 83 91 
<< m1 >>
rect 82 90 83 91 
<< m2 >>
rect 82 90 83 91 
<< m1 >>
rect 85 90 86 91 
<< m1 >>
rect 88 90 89 91 
<< m2 >>
rect 91 90 92 91 
<< m1 >>
rect 100 90 101 91 
<< m2 >>
rect 100 90 101 91 
<< m1 >>
rect 109 90 110 91 
<< m1 >>
rect 127 90 128 91 
<< m1 >>
rect 139 90 140 91 
<< m1 >>
rect 142 90 143 91 
<< m1 >>
rect 145 90 146 91 
<< m1 >>
rect 10 91 11 92 
<< m1 >>
rect 11 91 12 92 
<< m1 >>
rect 12 91 13 92 
<< m1 >>
rect 13 91 14 92 
<< m1 >>
rect 16 91 17 92 
<< m1 >>
rect 17 91 18 92 
<< m1 >>
rect 18 91 19 92 
<< m1 >>
rect 19 91 20 92 
<< m1 >>
rect 20 91 21 92 
<< m1 >>
rect 21 91 22 92 
<< m1 >>
rect 22 91 23 92 
<< m1 >>
rect 23 91 24 92 
<< m1 >>
rect 24 91 25 92 
<< m1 >>
rect 25 91 26 92 
<< m1 >>
rect 26 91 27 92 
<< m1 >>
rect 27 91 28 92 
<< m2 >>
rect 27 91 28 92 
<< m1 >>
rect 28 91 29 92 
<< m1 >>
rect 34 91 35 92 
<< m1 >>
rect 35 91 36 92 
<< m2 >>
rect 35 91 36 92 
<< m2c >>
rect 35 91 36 92 
<< m1 >>
rect 35 91 36 92 
<< m2 >>
rect 35 91 36 92 
<< m2 >>
rect 36 91 37 92 
<< m1 >>
rect 37 91 38 92 
<< m2 >>
rect 37 91 38 92 
<< m2 >>
rect 39 91 40 92 
<< m1 >>
rect 40 91 41 92 
<< m2 >>
rect 45 91 46 92 
<< m1 >>
rect 46 91 47 92 
<< m1 >>
rect 49 91 50 92 
<< m1 >>
rect 52 91 53 92 
<< m2 >>
rect 53 91 54 92 
<< m1 >>
rect 54 91 55 92 
<< m2 >>
rect 54 91 55 92 
<< m2c >>
rect 54 91 55 92 
<< m1 >>
rect 54 91 55 92 
<< m2 >>
rect 54 91 55 92 
<< m1 >>
rect 55 91 56 92 
<< m1 >>
rect 60 91 61 92 
<< m2 >>
rect 63 91 64 92 
<< m1 >>
rect 64 91 65 92 
<< m1 >>
rect 67 91 68 92 
<< m2 >>
rect 70 91 71 92 
<< m2 >>
rect 82 91 83 92 
<< m1 >>
rect 85 91 86 92 
<< m1 >>
rect 88 91 89 92 
<< m1 >>
rect 89 91 90 92 
<< m1 >>
rect 90 91 91 92 
<< m1 >>
rect 91 91 92 92 
<< m2 >>
rect 91 91 92 92 
<< m1 >>
rect 92 91 93 92 
<< m1 >>
rect 93 91 94 92 
<< m1 >>
rect 94 91 95 92 
<< m1 >>
rect 95 91 96 92 
<< m1 >>
rect 96 91 97 92 
<< m1 >>
rect 97 91 98 92 
<< m1 >>
rect 98 91 99 92 
<< m1 >>
rect 99 91 100 92 
<< m1 >>
rect 100 91 101 92 
<< m2 >>
rect 100 91 101 92 
<< m1 >>
rect 109 91 110 92 
<< m1 >>
rect 127 91 128 92 
<< m1 >>
rect 139 91 140 92 
<< m1 >>
rect 142 91 143 92 
<< m1 >>
rect 145 91 146 92 
<< m2 >>
rect 15 92 16 93 
<< m2 >>
rect 16 92 17 93 
<< m2 >>
rect 17 92 18 93 
<< m2 >>
rect 18 92 19 93 
<< m2 >>
rect 19 92 20 93 
<< m2 >>
rect 20 92 21 93 
<< m2 >>
rect 21 92 22 93 
<< m2 >>
rect 22 92 23 93 
<< m2 >>
rect 23 92 24 93 
<< m2 >>
rect 24 92 25 93 
<< m2 >>
rect 25 92 26 93 
<< m2 >>
rect 26 92 27 93 
<< m2 >>
rect 27 92 28 93 
<< m1 >>
rect 37 92 38 93 
<< m2 >>
rect 39 92 40 93 
<< m1 >>
rect 40 92 41 93 
<< m2 >>
rect 45 92 46 93 
<< m1 >>
rect 46 92 47 93 
<< m1 >>
rect 49 92 50 93 
<< m1 >>
rect 50 92 51 93 
<< m2 >>
rect 50 92 51 93 
<< m2c >>
rect 50 92 51 93 
<< m1 >>
rect 50 92 51 93 
<< m2 >>
rect 50 92 51 93 
<< m2 >>
rect 51 92 52 93 
<< m1 >>
rect 52 92 53 93 
<< m2 >>
rect 52 92 53 93 
<< m2 >>
rect 53 92 54 93 
<< m1 >>
rect 60 92 61 93 
<< m2 >>
rect 63 92 64 93 
<< m1 >>
rect 64 92 65 93 
<< m1 >>
rect 67 92 68 93 
<< m1 >>
rect 68 92 69 93 
<< m1 >>
rect 69 92 70 93 
<< m1 >>
rect 70 92 71 93 
<< m2 >>
rect 70 92 71 93 
<< m1 >>
rect 71 92 72 93 
<< m1 >>
rect 72 92 73 93 
<< m1 >>
rect 73 92 74 93 
<< m1 >>
rect 74 92 75 93 
<< m1 >>
rect 75 92 76 93 
<< m1 >>
rect 76 92 77 93 
<< m1 >>
rect 77 92 78 93 
<< m1 >>
rect 78 92 79 93 
<< m1 >>
rect 79 92 80 93 
<< m1 >>
rect 80 92 81 93 
<< m1 >>
rect 81 92 82 93 
<< m1 >>
rect 82 92 83 93 
<< m2 >>
rect 82 92 83 93 
<< m1 >>
rect 83 92 84 93 
<< m1 >>
rect 84 92 85 93 
<< m1 >>
rect 85 92 86 93 
<< m2 >>
rect 91 92 92 93 
<< m2 >>
rect 100 92 101 93 
<< m2 >>
rect 101 92 102 93 
<< m1 >>
rect 102 92 103 93 
<< m2 >>
rect 102 92 103 93 
<< m2c >>
rect 102 92 103 93 
<< m1 >>
rect 102 92 103 93 
<< m2 >>
rect 102 92 103 93 
<< m1 >>
rect 109 92 110 93 
<< m2 >>
rect 109 92 110 93 
<< m2c >>
rect 109 92 110 93 
<< m1 >>
rect 109 92 110 93 
<< m2 >>
rect 109 92 110 93 
<< m1 >>
rect 127 92 128 93 
<< m1 >>
rect 139 92 140 93 
<< m2 >>
rect 139 92 140 93 
<< m2c >>
rect 139 92 140 93 
<< m1 >>
rect 139 92 140 93 
<< m2 >>
rect 139 92 140 93 
<< m1 >>
rect 142 92 143 93 
<< m1 >>
rect 145 92 146 93 
<< m1 >>
rect 15 93 16 94 
<< m2 >>
rect 15 93 16 94 
<< m2c >>
rect 15 93 16 94 
<< m1 >>
rect 15 93 16 94 
<< m2 >>
rect 15 93 16 94 
<< m1 >>
rect 32 93 33 94 
<< m1 >>
rect 33 93 34 94 
<< m1 >>
rect 34 93 35 94 
<< m1 >>
rect 35 93 36 94 
<< m2 >>
rect 35 93 36 94 
<< m2c >>
rect 35 93 36 94 
<< m1 >>
rect 35 93 36 94 
<< m2 >>
rect 35 93 36 94 
<< m2 >>
rect 36 93 37 94 
<< m1 >>
rect 37 93 38 94 
<< m2 >>
rect 37 93 38 94 
<< m2 >>
rect 38 93 39 94 
<< m2 >>
rect 39 93 40 94 
<< m1 >>
rect 40 93 41 94 
<< m2 >>
rect 45 93 46 94 
<< m1 >>
rect 46 93 47 94 
<< m1 >>
rect 52 93 53 94 
<< m1 >>
rect 60 93 61 94 
<< m2 >>
rect 63 93 64 94 
<< m1 >>
rect 64 93 65 94 
<< m2 >>
rect 70 93 71 94 
<< m2 >>
rect 71 93 72 94 
<< m2 >>
rect 72 93 73 94 
<< m2 >>
rect 73 93 74 94 
<< m2 >>
rect 74 93 75 94 
<< m2 >>
rect 75 93 76 94 
<< m2 >>
rect 76 93 77 94 
<< m2 >>
rect 77 93 78 94 
<< m2 >>
rect 78 93 79 94 
<< m2 >>
rect 79 93 80 94 
<< m2 >>
rect 80 93 81 94 
<< m2 >>
rect 82 93 83 94 
<< m2 >>
rect 83 93 84 94 
<< m2 >>
rect 84 93 85 94 
<< m1 >>
rect 91 93 92 94 
<< m2 >>
rect 91 93 92 94 
<< m2c >>
rect 91 93 92 94 
<< m1 >>
rect 91 93 92 94 
<< m2 >>
rect 91 93 92 94 
<< m1 >>
rect 102 93 103 94 
<< m2 >>
rect 109 93 110 94 
<< m1 >>
rect 127 93 128 94 
<< m2 >>
rect 139 93 140 94 
<< m1 >>
rect 142 93 143 94 
<< m1 >>
rect 145 93 146 94 
<< m1 >>
rect 15 94 16 95 
<< m1 >>
rect 32 94 33 95 
<< m1 >>
rect 37 94 38 95 
<< m1 >>
rect 40 94 41 95 
<< m2 >>
rect 45 94 46 95 
<< m1 >>
rect 46 94 47 95 
<< m1 >>
rect 52 94 53 95 
<< m1 >>
rect 60 94 61 95 
<< m2 >>
rect 63 94 64 95 
<< m1 >>
rect 64 94 65 95 
<< m1 >>
rect 80 94 81 95 
<< m2 >>
rect 80 94 81 95 
<< m2c >>
rect 80 94 81 95 
<< m1 >>
rect 80 94 81 95 
<< m2 >>
rect 80 94 81 95 
<< m1 >>
rect 84 94 85 95 
<< m2 >>
rect 84 94 85 95 
<< m2c >>
rect 84 94 85 95 
<< m1 >>
rect 84 94 85 95 
<< m2 >>
rect 84 94 85 95 
<< m1 >>
rect 91 94 92 95 
<< m1 >>
rect 102 94 103 95 
<< m1 >>
rect 103 94 104 95 
<< m1 >>
rect 104 94 105 95 
<< m1 >>
rect 105 94 106 95 
<< m1 >>
rect 106 94 107 95 
<< m1 >>
rect 107 94 108 95 
<< m1 >>
rect 108 94 109 95 
<< m1 >>
rect 109 94 110 95 
<< m2 >>
rect 109 94 110 95 
<< m1 >>
rect 110 94 111 95 
<< m1 >>
rect 111 94 112 95 
<< m1 >>
rect 112 94 113 95 
<< m1 >>
rect 113 94 114 95 
<< m1 >>
rect 114 94 115 95 
<< m1 >>
rect 115 94 116 95 
<< m1 >>
rect 116 94 117 95 
<< m1 >>
rect 117 94 118 95 
<< m1 >>
rect 118 94 119 95 
<< m1 >>
rect 119 94 120 95 
<< m1 >>
rect 120 94 121 95 
<< m1 >>
rect 121 94 122 95 
<< m1 >>
rect 122 94 123 95 
<< m1 >>
rect 123 94 124 95 
<< m1 >>
rect 124 94 125 95 
<< m1 >>
rect 125 94 126 95 
<< m2 >>
rect 125 94 126 95 
<< m2c >>
rect 125 94 126 95 
<< m1 >>
rect 125 94 126 95 
<< m2 >>
rect 125 94 126 95 
<< m2 >>
rect 126 94 127 95 
<< m1 >>
rect 127 94 128 95 
<< m2 >>
rect 127 94 128 95 
<< m2 >>
rect 128 94 129 95 
<< m1 >>
rect 129 94 130 95 
<< m2 >>
rect 129 94 130 95 
<< m2c >>
rect 129 94 130 95 
<< m1 >>
rect 129 94 130 95 
<< m2 >>
rect 129 94 130 95 
<< m1 >>
rect 130 94 131 95 
<< m1 >>
rect 131 94 132 95 
<< m1 >>
rect 132 94 133 95 
<< m1 >>
rect 133 94 134 95 
<< m1 >>
rect 134 94 135 95 
<< m1 >>
rect 135 94 136 95 
<< m1 >>
rect 136 94 137 95 
<< m1 >>
rect 137 94 138 95 
<< m1 >>
rect 138 94 139 95 
<< m1 >>
rect 139 94 140 95 
<< m2 >>
rect 139 94 140 95 
<< m1 >>
rect 140 94 141 95 
<< m1 >>
rect 141 94 142 95 
<< m1 >>
rect 142 94 143 95 
<< m1 >>
rect 145 94 146 95 
<< m1 >>
rect 15 95 16 96 
<< m1 >>
rect 28 95 29 96 
<< m2 >>
rect 28 95 29 96 
<< m2c >>
rect 28 95 29 96 
<< m1 >>
rect 28 95 29 96 
<< m2 >>
rect 28 95 29 96 
<< m1 >>
rect 29 95 30 96 
<< m1 >>
rect 30 95 31 96 
<< m1 >>
rect 31 95 32 96 
<< m1 >>
rect 32 95 33 96 
<< m1 >>
rect 37 95 38 96 
<< m2 >>
rect 37 95 38 96 
<< m2c >>
rect 37 95 38 96 
<< m1 >>
rect 37 95 38 96 
<< m2 >>
rect 37 95 38 96 
<< m1 >>
rect 40 95 41 96 
<< m2 >>
rect 40 95 41 96 
<< m2c >>
rect 40 95 41 96 
<< m1 >>
rect 40 95 41 96 
<< m2 >>
rect 40 95 41 96 
<< m1 >>
rect 42 95 43 96 
<< m2 >>
rect 42 95 43 96 
<< m2c >>
rect 42 95 43 96 
<< m1 >>
rect 42 95 43 96 
<< m2 >>
rect 42 95 43 96 
<< m1 >>
rect 43 95 44 96 
<< m1 >>
rect 44 95 45 96 
<< m2 >>
rect 44 95 45 96 
<< m2c >>
rect 44 95 45 96 
<< m1 >>
rect 44 95 45 96 
<< m2 >>
rect 44 95 45 96 
<< m2 >>
rect 45 95 46 96 
<< m1 >>
rect 46 95 47 96 
<< m1 >>
rect 52 95 53 96 
<< m2 >>
rect 52 95 53 96 
<< m2c >>
rect 52 95 53 96 
<< m1 >>
rect 52 95 53 96 
<< m2 >>
rect 52 95 53 96 
<< m1 >>
rect 60 95 61 96 
<< m2 >>
rect 60 95 61 96 
<< m2c >>
rect 60 95 61 96 
<< m1 >>
rect 60 95 61 96 
<< m2 >>
rect 60 95 61 96 
<< m2 >>
rect 63 95 64 96 
<< m1 >>
rect 64 95 65 96 
<< m1 >>
rect 80 95 81 96 
<< m1 >>
rect 84 95 85 96 
<< m1 >>
rect 91 95 92 96 
<< m2 >>
rect 91 95 92 96 
<< m2c >>
rect 91 95 92 96 
<< m1 >>
rect 91 95 92 96 
<< m2 >>
rect 91 95 92 96 
<< m2 >>
rect 109 95 110 96 
<< m1 >>
rect 127 95 128 96 
<< m2 >>
rect 139 95 140 96 
<< m1 >>
rect 145 95 146 96 
<< m1 >>
rect 15 96 16 97 
<< m2 >>
rect 28 96 29 97 
<< m2 >>
rect 37 96 38 97 
<< m2 >>
rect 40 96 41 97 
<< m2 >>
rect 42 96 43 97 
<< m1 >>
rect 46 96 47 97 
<< m2 >>
rect 52 96 53 97 
<< m2 >>
rect 56 96 57 97 
<< m2 >>
rect 57 96 58 97 
<< m2 >>
rect 58 96 59 97 
<< m2 >>
rect 59 96 60 97 
<< m2 >>
rect 60 96 61 97 
<< m2 >>
rect 63 96 64 97 
<< m1 >>
rect 64 96 65 97 
<< m1 >>
rect 80 96 81 97 
<< m1 >>
rect 84 96 85 97 
<< m2 >>
rect 91 96 92 97 
<< m1 >>
rect 109 96 110 97 
<< m2 >>
rect 109 96 110 97 
<< m2c >>
rect 109 96 110 97 
<< m1 >>
rect 109 96 110 97 
<< m2 >>
rect 109 96 110 97 
<< m1 >>
rect 120 96 121 97 
<< m1 >>
rect 121 96 122 97 
<< m1 >>
rect 122 96 123 97 
<< m1 >>
rect 123 96 124 97 
<< m1 >>
rect 124 96 125 97 
<< m1 >>
rect 125 96 126 97 
<< m2 >>
rect 125 96 126 97 
<< m2c >>
rect 125 96 126 97 
<< m1 >>
rect 125 96 126 97 
<< m2 >>
rect 125 96 126 97 
<< m2 >>
rect 126 96 127 97 
<< m1 >>
rect 127 96 128 97 
<< m2 >>
rect 127 96 128 97 
<< m2 >>
rect 128 96 129 97 
<< m1 >>
rect 129 96 130 97 
<< m2 >>
rect 129 96 130 97 
<< m2c >>
rect 129 96 130 97 
<< m1 >>
rect 129 96 130 97 
<< m2 >>
rect 129 96 130 97 
<< m1 >>
rect 130 96 131 97 
<< m1 >>
rect 131 96 132 97 
<< m1 >>
rect 132 96 133 97 
<< m1 >>
rect 133 96 134 97 
<< m1 >>
rect 134 96 135 97 
<< m1 >>
rect 135 96 136 97 
<< m1 >>
rect 136 96 137 97 
<< m1 >>
rect 137 96 138 97 
<< m2 >>
rect 137 96 138 97 
<< m2c >>
rect 137 96 138 97 
<< m1 >>
rect 137 96 138 97 
<< m2 >>
rect 137 96 138 97 
<< m2 >>
rect 138 96 139 97 
<< m1 >>
rect 139 96 140 97 
<< m2 >>
rect 139 96 140 97 
<< m1 >>
rect 140 96 141 97 
<< m1 >>
rect 141 96 142 97 
<< m1 >>
rect 142 96 143 97 
<< m1 >>
rect 143 96 144 97 
<< m1 >>
rect 144 96 145 97 
<< m1 >>
rect 145 96 146 97 
<< m1 >>
rect 15 97 16 98 
<< m1 >>
rect 19 97 20 98 
<< m1 >>
rect 20 97 21 98 
<< m1 >>
rect 21 97 22 98 
<< m1 >>
rect 22 97 23 98 
<< m1 >>
rect 23 97 24 98 
<< m1 >>
rect 24 97 25 98 
<< m1 >>
rect 25 97 26 98 
<< m1 >>
rect 26 97 27 98 
<< m1 >>
rect 27 97 28 98 
<< m1 >>
rect 28 97 29 98 
<< m2 >>
rect 28 97 29 98 
<< m1 >>
rect 29 97 30 98 
<< m1 >>
rect 30 97 31 98 
<< m1 >>
rect 31 97 32 98 
<< m1 >>
rect 32 97 33 98 
<< m1 >>
rect 33 97 34 98 
<< m1 >>
rect 34 97 35 98 
<< m1 >>
rect 35 97 36 98 
<< m1 >>
rect 36 97 37 98 
<< m1 >>
rect 37 97 38 98 
<< m2 >>
rect 37 97 38 98 
<< m1 >>
rect 38 97 39 98 
<< m1 >>
rect 39 97 40 98 
<< m1 >>
rect 40 97 41 98 
<< m2 >>
rect 40 97 41 98 
<< m1 >>
rect 41 97 42 98 
<< m1 >>
rect 42 97 43 98 
<< m2 >>
rect 42 97 43 98 
<< m1 >>
rect 43 97 44 98 
<< m1 >>
rect 44 97 45 98 
<< m2 >>
rect 44 97 45 98 
<< m2c >>
rect 44 97 45 98 
<< m1 >>
rect 44 97 45 98 
<< m2 >>
rect 44 97 45 98 
<< m2 >>
rect 45 97 46 98 
<< m1 >>
rect 46 97 47 98 
<< m2 >>
rect 46 97 47 98 
<< m2 >>
rect 47 97 48 98 
<< m1 >>
rect 48 97 49 98 
<< m2 >>
rect 48 97 49 98 
<< m2c >>
rect 48 97 49 98 
<< m1 >>
rect 48 97 49 98 
<< m2 >>
rect 48 97 49 98 
<< m1 >>
rect 49 97 50 98 
<< m1 >>
rect 50 97 51 98 
<< m1 >>
rect 51 97 52 98 
<< m1 >>
rect 52 97 53 98 
<< m2 >>
rect 52 97 53 98 
<< m1 >>
rect 53 97 54 98 
<< m1 >>
rect 54 97 55 98 
<< m1 >>
rect 55 97 56 98 
<< m1 >>
rect 56 97 57 98 
<< m2 >>
rect 56 97 57 98 
<< m1 >>
rect 57 97 58 98 
<< m1 >>
rect 58 97 59 98 
<< m1 >>
rect 59 97 60 98 
<< m1 >>
rect 60 97 61 98 
<< m1 >>
rect 61 97 62 98 
<< m1 >>
rect 62 97 63 98 
<< m2 >>
rect 62 97 63 98 
<< m2c >>
rect 62 97 63 98 
<< m1 >>
rect 62 97 63 98 
<< m2 >>
rect 62 97 63 98 
<< m2 >>
rect 63 97 64 98 
<< m1 >>
rect 64 97 65 98 
<< m1 >>
rect 80 97 81 98 
<< m1 >>
rect 84 97 85 98 
<< m1 >>
rect 85 97 86 98 
<< m1 >>
rect 86 97 87 98 
<< m1 >>
rect 87 97 88 98 
<< m1 >>
rect 88 97 89 98 
<< m1 >>
rect 89 97 90 98 
<< m1 >>
rect 90 97 91 98 
<< m1 >>
rect 91 97 92 98 
<< m2 >>
rect 91 97 92 98 
<< m1 >>
rect 92 97 93 98 
<< m1 >>
rect 93 97 94 98 
<< m1 >>
rect 94 97 95 98 
<< m1 >>
rect 95 97 96 98 
<< m1 >>
rect 96 97 97 98 
<< m1 >>
rect 97 97 98 98 
<< m1 >>
rect 98 97 99 98 
<< m1 >>
rect 99 97 100 98 
<< m1 >>
rect 100 97 101 98 
<< m1 >>
rect 101 97 102 98 
<< m1 >>
rect 102 97 103 98 
<< m1 >>
rect 103 97 104 98 
<< m1 >>
rect 104 97 105 98 
<< m1 >>
rect 105 97 106 98 
<< m1 >>
rect 106 97 107 98 
<< m1 >>
rect 109 97 110 98 
<< m1 >>
rect 120 97 121 98 
<< m1 >>
rect 127 97 128 98 
<< m1 >>
rect 139 97 140 98 
<< m1 >>
rect 13 98 14 99 
<< m1 >>
rect 14 98 15 99 
<< m1 >>
rect 15 98 16 99 
<< m1 >>
rect 19 98 20 99 
<< m2 >>
rect 19 98 20 99 
<< m2c >>
rect 19 98 20 99 
<< m1 >>
rect 19 98 20 99 
<< m2 >>
rect 19 98 20 99 
<< m2 >>
rect 28 98 29 99 
<< m2 >>
rect 37 98 38 99 
<< m2 >>
rect 40 98 41 99 
<< m2 >>
rect 42 98 43 99 
<< m1 >>
rect 46 98 47 99 
<< m2 >>
rect 52 98 53 99 
<< m2 >>
rect 56 98 57 99 
<< m1 >>
rect 64 98 65 99 
<< m1 >>
rect 80 98 81 99 
<< m2 >>
rect 91 98 92 99 
<< m1 >>
rect 106 98 107 99 
<< m1 >>
rect 109 98 110 99 
<< m2 >>
rect 110 98 111 99 
<< m1 >>
rect 111 98 112 99 
<< m2 >>
rect 111 98 112 99 
<< m2c >>
rect 111 98 112 99 
<< m1 >>
rect 111 98 112 99 
<< m2 >>
rect 111 98 112 99 
<< m1 >>
rect 112 98 113 99 
<< m1 >>
rect 113 98 114 99 
<< m1 >>
rect 114 98 115 99 
<< m1 >>
rect 115 98 116 99 
<< m1 >>
rect 116 98 117 99 
<< m1 >>
rect 117 98 118 99 
<< m1 >>
rect 118 98 119 99 
<< m1 >>
rect 119 98 120 99 
<< m1 >>
rect 120 98 121 99 
<< m1 >>
rect 127 98 128 99 
<< m1 >>
rect 139 98 140 99 
<< m1 >>
rect 13 99 14 100 
<< m2 >>
rect 19 99 20 100 
<< m1 >>
rect 28 99 29 100 
<< m2 >>
rect 28 99 29 100 
<< m2c >>
rect 28 99 29 100 
<< m1 >>
rect 28 99 29 100 
<< m2 >>
rect 28 99 29 100 
<< m1 >>
rect 37 99 38 100 
<< m2 >>
rect 37 99 38 100 
<< m2c >>
rect 37 99 38 100 
<< m1 >>
rect 37 99 38 100 
<< m2 >>
rect 37 99 38 100 
<< m1 >>
rect 40 99 41 100 
<< m2 >>
rect 40 99 41 100 
<< m2c >>
rect 40 99 41 100 
<< m1 >>
rect 40 99 41 100 
<< m2 >>
rect 40 99 41 100 
<< m1 >>
rect 42 99 43 100 
<< m2 >>
rect 42 99 43 100 
<< m2c >>
rect 42 99 43 100 
<< m1 >>
rect 42 99 43 100 
<< m2 >>
rect 42 99 43 100 
<< m1 >>
rect 46 99 47 100 
<< m1 >>
rect 52 99 53 100 
<< m2 >>
rect 52 99 53 100 
<< m2c >>
rect 52 99 53 100 
<< m1 >>
rect 52 99 53 100 
<< m2 >>
rect 52 99 53 100 
<< m1 >>
rect 53 99 54 100 
<< m1 >>
rect 54 99 55 100 
<< m1 >>
rect 55 99 56 100 
<< m2 >>
rect 56 99 57 100 
<< m1 >>
rect 64 99 65 100 
<< m1 >>
rect 80 99 81 100 
<< m1 >>
rect 91 99 92 100 
<< m2 >>
rect 91 99 92 100 
<< m2c >>
rect 91 99 92 100 
<< m1 >>
rect 91 99 92 100 
<< m2 >>
rect 91 99 92 100 
<< m1 >>
rect 92 99 93 100 
<< m1 >>
rect 93 99 94 100 
<< m1 >>
rect 94 99 95 100 
<< m1 >>
rect 95 99 96 100 
<< m1 >>
rect 96 99 97 100 
<< m1 >>
rect 97 99 98 100 
<< m1 >>
rect 98 99 99 100 
<< m1 >>
rect 99 99 100 100 
<< m1 >>
rect 100 99 101 100 
<< m1 >>
rect 101 99 102 100 
<< m1 >>
rect 102 99 103 100 
<< m1 >>
rect 103 99 104 100 
<< m1 >>
rect 106 99 107 100 
<< m1 >>
rect 109 99 110 100 
<< m2 >>
rect 110 99 111 100 
<< m1 >>
rect 127 99 128 100 
<< m1 >>
rect 139 99 140 100 
<< m1 >>
rect 13 100 14 101 
<< m1 >>
rect 16 100 17 101 
<< m1 >>
rect 17 100 18 101 
<< m1 >>
rect 18 100 19 101 
<< m1 >>
rect 19 100 20 101 
<< m2 >>
rect 19 100 20 101 
<< m1 >>
rect 28 100 29 101 
<< m1 >>
rect 37 100 38 101 
<< m1 >>
rect 40 100 41 101 
<< m1 >>
rect 42 100 43 101 
<< m1 >>
rect 44 100 45 101 
<< m2 >>
rect 44 100 45 101 
<< m2c >>
rect 44 100 45 101 
<< m1 >>
rect 44 100 45 101 
<< m2 >>
rect 44 100 45 101 
<< m2 >>
rect 45 100 46 101 
<< m1 >>
rect 46 100 47 101 
<< m2 >>
rect 46 100 47 101 
<< m2 >>
rect 47 100 48 101 
<< m1 >>
rect 48 100 49 101 
<< m2 >>
rect 48 100 49 101 
<< m2c >>
rect 48 100 49 101 
<< m1 >>
rect 48 100 49 101 
<< m2 >>
rect 48 100 49 101 
<< m1 >>
rect 49 100 50 101 
<< m1 >>
rect 55 100 56 101 
<< m2 >>
rect 56 100 57 101 
<< m1 >>
rect 64 100 65 101 
<< m1 >>
rect 65 100 66 101 
<< m1 >>
rect 66 100 67 101 
<< m1 >>
rect 67 100 68 101 
<< m1 >>
rect 80 100 81 101 
<< m1 >>
rect 103 100 104 101 
<< m1 >>
rect 106 100 107 101 
<< m1 >>
rect 109 100 110 101 
<< m2 >>
rect 110 100 111 101 
<< m1 >>
rect 127 100 128 101 
<< m1 >>
rect 139 100 140 101 
<< m1 >>
rect 13 101 14 102 
<< m1 >>
rect 16 101 17 102 
<< m1 >>
rect 19 101 20 102 
<< m2 >>
rect 19 101 20 102 
<< m1 >>
rect 28 101 29 102 
<< m1 >>
rect 37 101 38 102 
<< m1 >>
rect 40 101 41 102 
<< m2 >>
rect 40 101 41 102 
<< m2c >>
rect 40 101 41 102 
<< m1 >>
rect 40 101 41 102 
<< m2 >>
rect 40 101 41 102 
<< m2 >>
rect 41 101 42 102 
<< m1 >>
rect 42 101 43 102 
<< m2 >>
rect 42 101 43 102 
<< m2 >>
rect 43 101 44 102 
<< m1 >>
rect 44 101 45 102 
<< m2 >>
rect 44 101 45 102 
<< m1 >>
rect 46 101 47 102 
<< m1 >>
rect 49 101 50 102 
<< m1 >>
rect 55 101 56 102 
<< m2 >>
rect 56 101 57 102 
<< m1 >>
rect 67 101 68 102 
<< m1 >>
rect 80 101 81 102 
<< m1 >>
rect 103 101 104 102 
<< m1 >>
rect 106 101 107 102 
<< m1 >>
rect 109 101 110 102 
<< m2 >>
rect 110 101 111 102 
<< m1 >>
rect 127 101 128 102 
<< m1 >>
rect 139 101 140 102 
<< pdiffusion >>
rect 12 102 13 103 
<< m1 >>
rect 13 102 14 103 
<< pdiffusion >>
rect 13 102 14 103 
<< pdiffusion >>
rect 14 102 15 103 
<< pdiffusion >>
rect 15 102 16 103 
<< m1 >>
rect 16 102 17 103 
<< pdiffusion >>
rect 16 102 17 103 
<< pdiffusion >>
rect 17 102 18 103 
<< m1 >>
rect 19 102 20 103 
<< m2 >>
rect 19 102 20 103 
<< m1 >>
rect 28 102 29 103 
<< pdiffusion >>
rect 30 102 31 103 
<< pdiffusion >>
rect 31 102 32 103 
<< pdiffusion >>
rect 32 102 33 103 
<< pdiffusion >>
rect 33 102 34 103 
<< pdiffusion >>
rect 34 102 35 103 
<< pdiffusion >>
rect 35 102 36 103 
<< m1 >>
rect 37 102 38 103 
<< m1 >>
rect 42 102 43 103 
<< m1 >>
rect 46 102 47 103 
<< pdiffusion >>
rect 48 102 49 103 
<< m1 >>
rect 49 102 50 103 
<< pdiffusion >>
rect 49 102 50 103 
<< pdiffusion >>
rect 50 102 51 103 
<< pdiffusion >>
rect 51 102 52 103 
<< pdiffusion >>
rect 52 102 53 103 
<< pdiffusion >>
rect 53 102 54 103 
<< m1 >>
rect 55 102 56 103 
<< m2 >>
rect 56 102 57 103 
<< pdiffusion >>
rect 66 102 67 103 
<< m1 >>
rect 67 102 68 103 
<< pdiffusion >>
rect 67 102 68 103 
<< pdiffusion >>
rect 68 102 69 103 
<< pdiffusion >>
rect 69 102 70 103 
<< pdiffusion >>
rect 70 102 71 103 
<< pdiffusion >>
rect 71 102 72 103 
<< m1 >>
rect 80 102 81 103 
<< pdiffusion >>
rect 84 102 85 103 
<< pdiffusion >>
rect 85 102 86 103 
<< pdiffusion >>
rect 86 102 87 103 
<< pdiffusion >>
rect 87 102 88 103 
<< pdiffusion >>
rect 88 102 89 103 
<< pdiffusion >>
rect 89 102 90 103 
<< pdiffusion >>
rect 102 102 103 103 
<< m1 >>
rect 103 102 104 103 
<< pdiffusion >>
rect 103 102 104 103 
<< pdiffusion >>
rect 104 102 105 103 
<< pdiffusion >>
rect 105 102 106 103 
<< m1 >>
rect 106 102 107 103 
<< pdiffusion >>
rect 106 102 107 103 
<< pdiffusion >>
rect 107 102 108 103 
<< m1 >>
rect 109 102 110 103 
<< m2 >>
rect 110 102 111 103 
<< pdiffusion >>
rect 120 102 121 103 
<< pdiffusion >>
rect 121 102 122 103 
<< pdiffusion >>
rect 122 102 123 103 
<< pdiffusion >>
rect 123 102 124 103 
<< pdiffusion >>
rect 124 102 125 103 
<< pdiffusion >>
rect 125 102 126 103 
<< m1 >>
rect 127 102 128 103 
<< pdiffusion >>
rect 138 102 139 103 
<< m1 >>
rect 139 102 140 103 
<< pdiffusion >>
rect 139 102 140 103 
<< pdiffusion >>
rect 140 102 141 103 
<< pdiffusion >>
rect 141 102 142 103 
<< pdiffusion >>
rect 142 102 143 103 
<< pdiffusion >>
rect 143 102 144 103 
<< pdiffusion >>
rect 12 103 13 104 
<< pdiffusion >>
rect 13 103 14 104 
<< pdiffusion >>
rect 14 103 15 104 
<< pdiffusion >>
rect 15 103 16 104 
<< pdiffusion >>
rect 16 103 17 104 
<< pdiffusion >>
rect 17 103 18 104 
<< m1 >>
rect 19 103 20 104 
<< m2 >>
rect 19 103 20 104 
<< m1 >>
rect 28 103 29 104 
<< pdiffusion >>
rect 30 103 31 104 
<< pdiffusion >>
rect 31 103 32 104 
<< pdiffusion >>
rect 32 103 33 104 
<< pdiffusion >>
rect 33 103 34 104 
<< pdiffusion >>
rect 34 103 35 104 
<< pdiffusion >>
rect 35 103 36 104 
<< m1 >>
rect 37 103 38 104 
<< m1 >>
rect 42 103 43 104 
<< m1 >>
rect 46 103 47 104 
<< pdiffusion >>
rect 48 103 49 104 
<< pdiffusion >>
rect 49 103 50 104 
<< pdiffusion >>
rect 50 103 51 104 
<< pdiffusion >>
rect 51 103 52 104 
<< pdiffusion >>
rect 52 103 53 104 
<< pdiffusion >>
rect 53 103 54 104 
<< m1 >>
rect 55 103 56 104 
<< m2 >>
rect 56 103 57 104 
<< pdiffusion >>
rect 66 103 67 104 
<< pdiffusion >>
rect 67 103 68 104 
<< pdiffusion >>
rect 68 103 69 104 
<< pdiffusion >>
rect 69 103 70 104 
<< pdiffusion >>
rect 70 103 71 104 
<< pdiffusion >>
rect 71 103 72 104 
<< m1 >>
rect 80 103 81 104 
<< pdiffusion >>
rect 84 103 85 104 
<< pdiffusion >>
rect 85 103 86 104 
<< pdiffusion >>
rect 86 103 87 104 
<< pdiffusion >>
rect 87 103 88 104 
<< pdiffusion >>
rect 88 103 89 104 
<< pdiffusion >>
rect 89 103 90 104 
<< pdiffusion >>
rect 102 103 103 104 
<< pdiffusion >>
rect 103 103 104 104 
<< pdiffusion >>
rect 104 103 105 104 
<< pdiffusion >>
rect 105 103 106 104 
<< pdiffusion >>
rect 106 103 107 104 
<< pdiffusion >>
rect 107 103 108 104 
<< m1 >>
rect 109 103 110 104 
<< m2 >>
rect 110 103 111 104 
<< pdiffusion >>
rect 120 103 121 104 
<< pdiffusion >>
rect 121 103 122 104 
<< pdiffusion >>
rect 122 103 123 104 
<< pdiffusion >>
rect 123 103 124 104 
<< pdiffusion >>
rect 124 103 125 104 
<< pdiffusion >>
rect 125 103 126 104 
<< m1 >>
rect 127 103 128 104 
<< pdiffusion >>
rect 138 103 139 104 
<< pdiffusion >>
rect 139 103 140 104 
<< pdiffusion >>
rect 140 103 141 104 
<< pdiffusion >>
rect 141 103 142 104 
<< pdiffusion >>
rect 142 103 143 104 
<< pdiffusion >>
rect 143 103 144 104 
<< pdiffusion >>
rect 12 104 13 105 
<< pdiffusion >>
rect 13 104 14 105 
<< pdiffusion >>
rect 14 104 15 105 
<< pdiffusion >>
rect 15 104 16 105 
<< pdiffusion >>
rect 16 104 17 105 
<< pdiffusion >>
rect 17 104 18 105 
<< m1 >>
rect 19 104 20 105 
<< m2 >>
rect 19 104 20 105 
<< m1 >>
rect 28 104 29 105 
<< pdiffusion >>
rect 30 104 31 105 
<< pdiffusion >>
rect 31 104 32 105 
<< pdiffusion >>
rect 32 104 33 105 
<< pdiffusion >>
rect 33 104 34 105 
<< pdiffusion >>
rect 34 104 35 105 
<< pdiffusion >>
rect 35 104 36 105 
<< m1 >>
rect 37 104 38 105 
<< m1 >>
rect 42 104 43 105 
<< m1 >>
rect 46 104 47 105 
<< pdiffusion >>
rect 48 104 49 105 
<< pdiffusion >>
rect 49 104 50 105 
<< pdiffusion >>
rect 50 104 51 105 
<< pdiffusion >>
rect 51 104 52 105 
<< pdiffusion >>
rect 52 104 53 105 
<< pdiffusion >>
rect 53 104 54 105 
<< m1 >>
rect 55 104 56 105 
<< m2 >>
rect 56 104 57 105 
<< pdiffusion >>
rect 66 104 67 105 
<< pdiffusion >>
rect 67 104 68 105 
<< pdiffusion >>
rect 68 104 69 105 
<< pdiffusion >>
rect 69 104 70 105 
<< pdiffusion >>
rect 70 104 71 105 
<< pdiffusion >>
rect 71 104 72 105 
<< m1 >>
rect 80 104 81 105 
<< pdiffusion >>
rect 84 104 85 105 
<< pdiffusion >>
rect 85 104 86 105 
<< pdiffusion >>
rect 86 104 87 105 
<< pdiffusion >>
rect 87 104 88 105 
<< pdiffusion >>
rect 88 104 89 105 
<< pdiffusion >>
rect 89 104 90 105 
<< pdiffusion >>
rect 102 104 103 105 
<< pdiffusion >>
rect 103 104 104 105 
<< pdiffusion >>
rect 104 104 105 105 
<< pdiffusion >>
rect 105 104 106 105 
<< pdiffusion >>
rect 106 104 107 105 
<< pdiffusion >>
rect 107 104 108 105 
<< m1 >>
rect 109 104 110 105 
<< m2 >>
rect 110 104 111 105 
<< pdiffusion >>
rect 120 104 121 105 
<< pdiffusion >>
rect 121 104 122 105 
<< pdiffusion >>
rect 122 104 123 105 
<< pdiffusion >>
rect 123 104 124 105 
<< pdiffusion >>
rect 124 104 125 105 
<< pdiffusion >>
rect 125 104 126 105 
<< m1 >>
rect 127 104 128 105 
<< pdiffusion >>
rect 138 104 139 105 
<< pdiffusion >>
rect 139 104 140 105 
<< pdiffusion >>
rect 140 104 141 105 
<< pdiffusion >>
rect 141 104 142 105 
<< pdiffusion >>
rect 142 104 143 105 
<< pdiffusion >>
rect 143 104 144 105 
<< pdiffusion >>
rect 12 105 13 106 
<< pdiffusion >>
rect 13 105 14 106 
<< pdiffusion >>
rect 14 105 15 106 
<< pdiffusion >>
rect 15 105 16 106 
<< pdiffusion >>
rect 16 105 17 106 
<< pdiffusion >>
rect 17 105 18 106 
<< m1 >>
rect 19 105 20 106 
<< m2 >>
rect 19 105 20 106 
<< m1 >>
rect 28 105 29 106 
<< pdiffusion >>
rect 30 105 31 106 
<< pdiffusion >>
rect 31 105 32 106 
<< pdiffusion >>
rect 32 105 33 106 
<< pdiffusion >>
rect 33 105 34 106 
<< pdiffusion >>
rect 34 105 35 106 
<< pdiffusion >>
rect 35 105 36 106 
<< m1 >>
rect 37 105 38 106 
<< m1 >>
rect 42 105 43 106 
<< m1 >>
rect 46 105 47 106 
<< pdiffusion >>
rect 48 105 49 106 
<< pdiffusion >>
rect 49 105 50 106 
<< pdiffusion >>
rect 50 105 51 106 
<< pdiffusion >>
rect 51 105 52 106 
<< pdiffusion >>
rect 52 105 53 106 
<< pdiffusion >>
rect 53 105 54 106 
<< m1 >>
rect 55 105 56 106 
<< m2 >>
rect 56 105 57 106 
<< pdiffusion >>
rect 66 105 67 106 
<< pdiffusion >>
rect 67 105 68 106 
<< pdiffusion >>
rect 68 105 69 106 
<< pdiffusion >>
rect 69 105 70 106 
<< pdiffusion >>
rect 70 105 71 106 
<< pdiffusion >>
rect 71 105 72 106 
<< m1 >>
rect 80 105 81 106 
<< pdiffusion >>
rect 84 105 85 106 
<< pdiffusion >>
rect 85 105 86 106 
<< pdiffusion >>
rect 86 105 87 106 
<< pdiffusion >>
rect 87 105 88 106 
<< pdiffusion >>
rect 88 105 89 106 
<< pdiffusion >>
rect 89 105 90 106 
<< pdiffusion >>
rect 102 105 103 106 
<< pdiffusion >>
rect 103 105 104 106 
<< pdiffusion >>
rect 104 105 105 106 
<< pdiffusion >>
rect 105 105 106 106 
<< pdiffusion >>
rect 106 105 107 106 
<< pdiffusion >>
rect 107 105 108 106 
<< m1 >>
rect 109 105 110 106 
<< m2 >>
rect 110 105 111 106 
<< pdiffusion >>
rect 120 105 121 106 
<< pdiffusion >>
rect 121 105 122 106 
<< pdiffusion >>
rect 122 105 123 106 
<< pdiffusion >>
rect 123 105 124 106 
<< pdiffusion >>
rect 124 105 125 106 
<< pdiffusion >>
rect 125 105 126 106 
<< m1 >>
rect 127 105 128 106 
<< pdiffusion >>
rect 138 105 139 106 
<< pdiffusion >>
rect 139 105 140 106 
<< pdiffusion >>
rect 140 105 141 106 
<< pdiffusion >>
rect 141 105 142 106 
<< pdiffusion >>
rect 142 105 143 106 
<< pdiffusion >>
rect 143 105 144 106 
<< pdiffusion >>
rect 12 106 13 107 
<< pdiffusion >>
rect 13 106 14 107 
<< pdiffusion >>
rect 14 106 15 107 
<< pdiffusion >>
rect 15 106 16 107 
<< pdiffusion >>
rect 16 106 17 107 
<< pdiffusion >>
rect 17 106 18 107 
<< m1 >>
rect 19 106 20 107 
<< m2 >>
rect 19 106 20 107 
<< m1 >>
rect 28 106 29 107 
<< pdiffusion >>
rect 30 106 31 107 
<< pdiffusion >>
rect 31 106 32 107 
<< pdiffusion >>
rect 32 106 33 107 
<< pdiffusion >>
rect 33 106 34 107 
<< pdiffusion >>
rect 34 106 35 107 
<< pdiffusion >>
rect 35 106 36 107 
<< m1 >>
rect 37 106 38 107 
<< m1 >>
rect 42 106 43 107 
<< m1 >>
rect 46 106 47 107 
<< pdiffusion >>
rect 48 106 49 107 
<< pdiffusion >>
rect 49 106 50 107 
<< pdiffusion >>
rect 50 106 51 107 
<< pdiffusion >>
rect 51 106 52 107 
<< pdiffusion >>
rect 52 106 53 107 
<< pdiffusion >>
rect 53 106 54 107 
<< m1 >>
rect 55 106 56 107 
<< m2 >>
rect 56 106 57 107 
<< pdiffusion >>
rect 66 106 67 107 
<< pdiffusion >>
rect 67 106 68 107 
<< pdiffusion >>
rect 68 106 69 107 
<< pdiffusion >>
rect 69 106 70 107 
<< pdiffusion >>
rect 70 106 71 107 
<< pdiffusion >>
rect 71 106 72 107 
<< m1 >>
rect 80 106 81 107 
<< pdiffusion >>
rect 84 106 85 107 
<< pdiffusion >>
rect 85 106 86 107 
<< pdiffusion >>
rect 86 106 87 107 
<< pdiffusion >>
rect 87 106 88 107 
<< pdiffusion >>
rect 88 106 89 107 
<< pdiffusion >>
rect 89 106 90 107 
<< pdiffusion >>
rect 102 106 103 107 
<< pdiffusion >>
rect 103 106 104 107 
<< pdiffusion >>
rect 104 106 105 107 
<< pdiffusion >>
rect 105 106 106 107 
<< pdiffusion >>
rect 106 106 107 107 
<< pdiffusion >>
rect 107 106 108 107 
<< m1 >>
rect 109 106 110 107 
<< m2 >>
rect 110 106 111 107 
<< pdiffusion >>
rect 120 106 121 107 
<< pdiffusion >>
rect 121 106 122 107 
<< pdiffusion >>
rect 122 106 123 107 
<< pdiffusion >>
rect 123 106 124 107 
<< pdiffusion >>
rect 124 106 125 107 
<< pdiffusion >>
rect 125 106 126 107 
<< m1 >>
rect 127 106 128 107 
<< pdiffusion >>
rect 138 106 139 107 
<< pdiffusion >>
rect 139 106 140 107 
<< pdiffusion >>
rect 140 106 141 107 
<< pdiffusion >>
rect 141 106 142 107 
<< pdiffusion >>
rect 142 106 143 107 
<< pdiffusion >>
rect 143 106 144 107 
<< pdiffusion >>
rect 12 107 13 108 
<< m1 >>
rect 13 107 14 108 
<< pdiffusion >>
rect 13 107 14 108 
<< pdiffusion >>
rect 14 107 15 108 
<< pdiffusion >>
rect 15 107 16 108 
<< pdiffusion >>
rect 16 107 17 108 
<< pdiffusion >>
rect 17 107 18 108 
<< m1 >>
rect 19 107 20 108 
<< m2 >>
rect 19 107 20 108 
<< m1 >>
rect 28 107 29 108 
<< pdiffusion >>
rect 30 107 31 108 
<< pdiffusion >>
rect 31 107 32 108 
<< pdiffusion >>
rect 32 107 33 108 
<< pdiffusion >>
rect 33 107 34 108 
<< pdiffusion >>
rect 34 107 35 108 
<< pdiffusion >>
rect 35 107 36 108 
<< m1 >>
rect 37 107 38 108 
<< m1 >>
rect 42 107 43 108 
<< m1 >>
rect 46 107 47 108 
<< pdiffusion >>
rect 48 107 49 108 
<< m1 >>
rect 49 107 50 108 
<< pdiffusion >>
rect 49 107 50 108 
<< pdiffusion >>
rect 50 107 51 108 
<< pdiffusion >>
rect 51 107 52 108 
<< pdiffusion >>
rect 52 107 53 108 
<< pdiffusion >>
rect 53 107 54 108 
<< m1 >>
rect 55 107 56 108 
<< m2 >>
rect 56 107 57 108 
<< pdiffusion >>
rect 66 107 67 108 
<< pdiffusion >>
rect 67 107 68 108 
<< pdiffusion >>
rect 68 107 69 108 
<< pdiffusion >>
rect 69 107 70 108 
<< pdiffusion >>
rect 70 107 71 108 
<< pdiffusion >>
rect 71 107 72 108 
<< m1 >>
rect 80 107 81 108 
<< pdiffusion >>
rect 84 107 85 108 
<< m1 >>
rect 85 107 86 108 
<< pdiffusion >>
rect 85 107 86 108 
<< pdiffusion >>
rect 86 107 87 108 
<< pdiffusion >>
rect 87 107 88 108 
<< m1 >>
rect 88 107 89 108 
<< pdiffusion >>
rect 88 107 89 108 
<< pdiffusion >>
rect 89 107 90 108 
<< pdiffusion >>
rect 102 107 103 108 
<< pdiffusion >>
rect 103 107 104 108 
<< pdiffusion >>
rect 104 107 105 108 
<< pdiffusion >>
rect 105 107 106 108 
<< pdiffusion >>
rect 106 107 107 108 
<< pdiffusion >>
rect 107 107 108 108 
<< m1 >>
rect 109 107 110 108 
<< m2 >>
rect 110 107 111 108 
<< pdiffusion >>
rect 120 107 121 108 
<< pdiffusion >>
rect 121 107 122 108 
<< pdiffusion >>
rect 122 107 123 108 
<< pdiffusion >>
rect 123 107 124 108 
<< m1 >>
rect 124 107 125 108 
<< pdiffusion >>
rect 124 107 125 108 
<< pdiffusion >>
rect 125 107 126 108 
<< m1 >>
rect 127 107 128 108 
<< pdiffusion >>
rect 138 107 139 108 
<< pdiffusion >>
rect 139 107 140 108 
<< pdiffusion >>
rect 140 107 141 108 
<< pdiffusion >>
rect 141 107 142 108 
<< pdiffusion >>
rect 142 107 143 108 
<< pdiffusion >>
rect 143 107 144 108 
<< m1 >>
rect 13 108 14 109 
<< m1 >>
rect 19 108 20 109 
<< m2 >>
rect 19 108 20 109 
<< m1 >>
rect 28 108 29 109 
<< m1 >>
rect 37 108 38 109 
<< m1 >>
rect 42 108 43 109 
<< m1 >>
rect 46 108 47 109 
<< m1 >>
rect 49 108 50 109 
<< m1 >>
rect 55 108 56 109 
<< m2 >>
rect 56 108 57 109 
<< m1 >>
rect 80 108 81 109 
<< m1 >>
rect 85 108 86 109 
<< m1 >>
rect 88 108 89 109 
<< m1 >>
rect 109 108 110 109 
<< m2 >>
rect 110 108 111 109 
<< m1 >>
rect 124 108 125 109 
<< m1 >>
rect 127 108 128 109 
<< m1 >>
rect 13 109 14 110 
<< m1 >>
rect 19 109 20 110 
<< m2 >>
rect 19 109 20 110 
<< m1 >>
rect 28 109 29 110 
<< m1 >>
rect 37 109 38 110 
<< m1 >>
rect 42 109 43 110 
<< m1 >>
rect 46 109 47 110 
<< m1 >>
rect 49 109 50 110 
<< m1 >>
rect 53 109 54 110 
<< m2 >>
rect 53 109 54 110 
<< m2c >>
rect 53 109 54 110 
<< m1 >>
rect 53 109 54 110 
<< m2 >>
rect 53 109 54 110 
<< m2 >>
rect 54 109 55 110 
<< m1 >>
rect 55 109 56 110 
<< m2 >>
rect 55 109 56 110 
<< m2 >>
rect 56 109 57 110 
<< m1 >>
rect 76 109 77 110 
<< m1 >>
rect 77 109 78 110 
<< m1 >>
rect 78 109 79 110 
<< m2 >>
rect 78 109 79 110 
<< m2c >>
rect 78 109 79 110 
<< m1 >>
rect 78 109 79 110 
<< m2 >>
rect 78 109 79 110 
<< m2 >>
rect 79 109 80 110 
<< m1 >>
rect 80 109 81 110 
<< m2 >>
rect 80 109 81 110 
<< m2 >>
rect 81 109 82 110 
<< m1 >>
rect 82 109 83 110 
<< m2 >>
rect 82 109 83 110 
<< m2c >>
rect 82 109 83 110 
<< m1 >>
rect 82 109 83 110 
<< m2 >>
rect 82 109 83 110 
<< m1 >>
rect 83 109 84 110 
<< m1 >>
rect 84 109 85 110 
<< m1 >>
rect 85 109 86 110 
<< m1 >>
rect 88 109 89 110 
<< m1 >>
rect 89 109 90 110 
<< m1 >>
rect 107 109 108 110 
<< m2 >>
rect 107 109 108 110 
<< m2c >>
rect 107 109 108 110 
<< m1 >>
rect 107 109 108 110 
<< m2 >>
rect 107 109 108 110 
<< m2 >>
rect 108 109 109 110 
<< m1 >>
rect 109 109 110 110 
<< m2 >>
rect 109 109 110 110 
<< m2 >>
rect 110 109 111 110 
<< m1 >>
rect 124 109 125 110 
<< m1 >>
rect 127 109 128 110 
<< m1 >>
rect 13 110 14 111 
<< m1 >>
rect 14 110 15 111 
<< m1 >>
rect 15 110 16 111 
<< m1 >>
rect 16 110 17 111 
<< m1 >>
rect 17 110 18 111 
<< m2 >>
rect 17 110 18 111 
<< m2c >>
rect 17 110 18 111 
<< m1 >>
rect 17 110 18 111 
<< m2 >>
rect 17 110 18 111 
<< m2 >>
rect 18 110 19 111 
<< m1 >>
rect 19 110 20 111 
<< m2 >>
rect 19 110 20 111 
<< m1 >>
rect 28 110 29 111 
<< m1 >>
rect 29 110 30 111 
<< m1 >>
rect 30 110 31 111 
<< m2 >>
rect 30 110 31 111 
<< m2c >>
rect 30 110 31 111 
<< m1 >>
rect 30 110 31 111 
<< m2 >>
rect 30 110 31 111 
<< m1 >>
rect 37 110 38 111 
<< m2 >>
rect 37 110 38 111 
<< m2c >>
rect 37 110 38 111 
<< m1 >>
rect 37 110 38 111 
<< m2 >>
rect 37 110 38 111 
<< m1 >>
rect 42 110 43 111 
<< m2 >>
rect 42 110 43 111 
<< m2c >>
rect 42 110 43 111 
<< m1 >>
rect 42 110 43 111 
<< m2 >>
rect 42 110 43 111 
<< m1 >>
rect 46 110 47 111 
<< m1 >>
rect 49 110 50 111 
<< m1 >>
rect 52 110 53 111 
<< m1 >>
rect 53 110 54 111 
<< m1 >>
rect 55 110 56 111 
<< m1 >>
rect 76 110 77 111 
<< m2 >>
rect 76 110 77 111 
<< m2c >>
rect 76 110 77 111 
<< m1 >>
rect 76 110 77 111 
<< m2 >>
rect 76 110 77 111 
<< m1 >>
rect 80 110 81 111 
<< m1 >>
rect 89 110 90 111 
<< m2 >>
rect 89 110 90 111 
<< m2c >>
rect 89 110 90 111 
<< m1 >>
rect 89 110 90 111 
<< m2 >>
rect 89 110 90 111 
<< m1 >>
rect 107 110 108 111 
<< m1 >>
rect 109 110 110 111 
<< m1 >>
rect 124 110 125 111 
<< m1 >>
rect 127 110 128 111 
<< m1 >>
rect 19 111 20 112 
<< m2 >>
rect 30 111 31 112 
<< m2 >>
rect 37 111 38 112 
<< m2 >>
rect 42 111 43 112 
<< m1 >>
rect 46 111 47 112 
<< m1 >>
rect 49 111 50 112 
<< m1 >>
rect 52 111 53 112 
<< m1 >>
rect 55 111 56 112 
<< m2 >>
rect 76 111 77 112 
<< m1 >>
rect 80 111 81 112 
<< m2 >>
rect 89 111 90 112 
<< m1 >>
rect 107 111 108 112 
<< m1 >>
rect 109 111 110 112 
<< m1 >>
rect 124 111 125 112 
<< m1 >>
rect 127 111 128 112 
<< m1 >>
rect 19 112 20 113 
<< m1 >>
rect 20 112 21 113 
<< m1 >>
rect 21 112 22 113 
<< m1 >>
rect 22 112 23 113 
<< m1 >>
rect 23 112 24 113 
<< m1 >>
rect 24 112 25 113 
<< m1 >>
rect 25 112 26 113 
<< m1 >>
rect 26 112 27 113 
<< m1 >>
rect 27 112 28 113 
<< m1 >>
rect 28 112 29 113 
<< m1 >>
rect 29 112 30 113 
<< m1 >>
rect 30 112 31 113 
<< m2 >>
rect 30 112 31 113 
<< m1 >>
rect 31 112 32 113 
<< m1 >>
rect 32 112 33 113 
<< m1 >>
rect 33 112 34 113 
<< m1 >>
rect 34 112 35 113 
<< m1 >>
rect 35 112 36 113 
<< m1 >>
rect 36 112 37 113 
<< m1 >>
rect 37 112 38 113 
<< m2 >>
rect 37 112 38 113 
<< m1 >>
rect 38 112 39 113 
<< m1 >>
rect 39 112 40 113 
<< m1 >>
rect 40 112 41 113 
<< m1 >>
rect 41 112 42 113 
<< m1 >>
rect 42 112 43 113 
<< m2 >>
rect 42 112 43 113 
<< m1 >>
rect 43 112 44 113 
<< m1 >>
rect 44 112 45 113 
<< m2 >>
rect 44 112 45 113 
<< m2c >>
rect 44 112 45 113 
<< m1 >>
rect 44 112 45 113 
<< m2 >>
rect 44 112 45 113 
<< m2 >>
rect 45 112 46 113 
<< m1 >>
rect 46 112 47 113 
<< m2 >>
rect 46 112 47 113 
<< m2 >>
rect 47 112 48 113 
<< m1 >>
rect 48 112 49 113 
<< m2 >>
rect 48 112 49 113 
<< m2c >>
rect 48 112 49 113 
<< m1 >>
rect 48 112 49 113 
<< m2 >>
rect 48 112 49 113 
<< m1 >>
rect 49 112 50 113 
<< m1 >>
rect 52 112 53 113 
<< m1 >>
rect 55 112 56 113 
<< m1 >>
rect 56 112 57 113 
<< m1 >>
rect 57 112 58 113 
<< m1 >>
rect 58 112 59 113 
<< m1 >>
rect 59 112 60 113 
<< m1 >>
rect 60 112 61 113 
<< m1 >>
rect 61 112 62 113 
<< m1 >>
rect 62 112 63 113 
<< m1 >>
rect 63 112 64 113 
<< m1 >>
rect 64 112 65 113 
<< m1 >>
rect 65 112 66 113 
<< m1 >>
rect 66 112 67 113 
<< m1 >>
rect 67 112 68 113 
<< m1 >>
rect 68 112 69 113 
<< m1 >>
rect 69 112 70 113 
<< m1 >>
rect 70 112 71 113 
<< m1 >>
rect 71 112 72 113 
<< m1 >>
rect 72 112 73 113 
<< m1 >>
rect 73 112 74 113 
<< m1 >>
rect 74 112 75 113 
<< m1 >>
rect 75 112 76 113 
<< m1 >>
rect 76 112 77 113 
<< m2 >>
rect 76 112 77 113 
<< m1 >>
rect 77 112 78 113 
<< m1 >>
rect 78 112 79 113 
<< m2 >>
rect 78 112 79 113 
<< m2c >>
rect 78 112 79 113 
<< m1 >>
rect 78 112 79 113 
<< m2 >>
rect 78 112 79 113 
<< m2 >>
rect 79 112 80 113 
<< m1 >>
rect 80 112 81 113 
<< m2 >>
rect 80 112 81 113 
<< m2 >>
rect 81 112 82 113 
<< m1 >>
rect 82 112 83 113 
<< m2 >>
rect 82 112 83 113 
<< m2c >>
rect 82 112 83 113 
<< m1 >>
rect 82 112 83 113 
<< m2 >>
rect 82 112 83 113 
<< m1 >>
rect 83 112 84 113 
<< m1 >>
rect 84 112 85 113 
<< m1 >>
rect 85 112 86 113 
<< m2 >>
rect 86 112 87 113 
<< m1 >>
rect 87 112 88 113 
<< m2 >>
rect 87 112 88 113 
<< m2c >>
rect 87 112 88 113 
<< m1 >>
rect 87 112 88 113 
<< m2 >>
rect 87 112 88 113 
<< m1 >>
rect 88 112 89 113 
<< m1 >>
rect 89 112 90 113 
<< m2 >>
rect 89 112 90 113 
<< m1 >>
rect 90 112 91 113 
<< m2 >>
rect 90 112 91 113 
<< m1 >>
rect 91 112 92 113 
<< m2 >>
rect 91 112 92 113 
<< m1 >>
rect 92 112 93 113 
<< m2 >>
rect 92 112 93 113 
<< m1 >>
rect 93 112 94 113 
<< m2 >>
rect 93 112 94 113 
<< m1 >>
rect 94 112 95 113 
<< m2 >>
rect 94 112 95 113 
<< m1 >>
rect 95 112 96 113 
<< m2 >>
rect 95 112 96 113 
<< m1 >>
rect 96 112 97 113 
<< m2 >>
rect 96 112 97 113 
<< m1 >>
rect 97 112 98 113 
<< m2 >>
rect 97 112 98 113 
<< m1 >>
rect 98 112 99 113 
<< m2 >>
rect 98 112 99 113 
<< m1 >>
rect 99 112 100 113 
<< m2 >>
rect 99 112 100 113 
<< m1 >>
rect 100 112 101 113 
<< m2 >>
rect 100 112 101 113 
<< m1 >>
rect 101 112 102 113 
<< m2 >>
rect 101 112 102 113 
<< m1 >>
rect 102 112 103 113 
<< m2 >>
rect 102 112 103 113 
<< m1 >>
rect 103 112 104 113 
<< m2 >>
rect 103 112 104 113 
<< m1 >>
rect 104 112 105 113 
<< m2 >>
rect 104 112 105 113 
<< m1 >>
rect 105 112 106 113 
<< m2 >>
rect 105 112 106 113 
<< m1 >>
rect 106 112 107 113 
<< m2 >>
rect 106 112 107 113 
<< m1 >>
rect 107 112 108 113 
<< m2 >>
rect 107 112 108 113 
<< m2 >>
rect 108 112 109 113 
<< m1 >>
rect 109 112 110 113 
<< m2 >>
rect 109 112 110 113 
<< m2 >>
rect 110 112 111 113 
<< m1 >>
rect 111 112 112 113 
<< m2 >>
rect 111 112 112 113 
<< m2c >>
rect 111 112 112 113 
<< m1 >>
rect 111 112 112 113 
<< m2 >>
rect 111 112 112 113 
<< m1 >>
rect 112 112 113 113 
<< m1 >>
rect 113 112 114 113 
<< m1 >>
rect 114 112 115 113 
<< m1 >>
rect 115 112 116 113 
<< m1 >>
rect 116 112 117 113 
<< m1 >>
rect 117 112 118 113 
<< m1 >>
rect 118 112 119 113 
<< m1 >>
rect 119 112 120 113 
<< m1 >>
rect 120 112 121 113 
<< m1 >>
rect 121 112 122 113 
<< m1 >>
rect 122 112 123 113 
<< m1 >>
rect 123 112 124 113 
<< m1 >>
rect 124 112 125 113 
<< m1 >>
rect 127 112 128 113 
<< m2 >>
rect 30 113 31 114 
<< m2 >>
rect 37 113 38 114 
<< m2 >>
rect 42 113 43 114 
<< m1 >>
rect 46 113 47 114 
<< m1 >>
rect 52 113 53 114 
<< m2 >>
rect 76 113 77 114 
<< m1 >>
rect 80 113 81 114 
<< m1 >>
rect 85 113 86 114 
<< m2 >>
rect 86 113 87 114 
<< m1 >>
rect 109 113 110 114 
<< m1 >>
rect 127 113 128 114 
<< m2 >>
rect 30 114 31 115 
<< m1 >>
rect 31 114 32 115 
<< m1 >>
rect 32 114 33 115 
<< m1 >>
rect 33 114 34 115 
<< m1 >>
rect 34 114 35 115 
<< m1 >>
rect 35 114 36 115 
<< m1 >>
rect 36 114 37 115 
<< m1 >>
rect 37 114 38 115 
<< m2 >>
rect 37 114 38 115 
<< m2c >>
rect 37 114 38 115 
<< m1 >>
rect 37 114 38 115 
<< m2 >>
rect 37 114 38 115 
<< m1 >>
rect 42 114 43 115 
<< m2 >>
rect 42 114 43 115 
<< m2c >>
rect 42 114 43 115 
<< m1 >>
rect 42 114 43 115 
<< m2 >>
rect 42 114 43 115 
<< m1 >>
rect 43 114 44 115 
<< m1 >>
rect 44 114 45 115 
<< m2 >>
rect 44 114 45 115 
<< m2c >>
rect 44 114 45 115 
<< m1 >>
rect 44 114 45 115 
<< m2 >>
rect 44 114 45 115 
<< m2 >>
rect 45 114 46 115 
<< m1 >>
rect 46 114 47 115 
<< m2 >>
rect 46 114 47 115 
<< m2 >>
rect 47 114 48 115 
<< m1 >>
rect 48 114 49 115 
<< m2 >>
rect 48 114 49 115 
<< m2c >>
rect 48 114 49 115 
<< m1 >>
rect 48 114 49 115 
<< m2 >>
rect 48 114 49 115 
<< m1 >>
rect 49 114 50 115 
<< m1 >>
rect 50 114 51 115 
<< m2 >>
rect 50 114 51 115 
<< m2c >>
rect 50 114 51 115 
<< m1 >>
rect 50 114 51 115 
<< m2 >>
rect 50 114 51 115 
<< m2 >>
rect 51 114 52 115 
<< m1 >>
rect 52 114 53 115 
<< m2 >>
rect 52 114 53 115 
<< m2 >>
rect 53 114 54 115 
<< m1 >>
rect 54 114 55 115 
<< m2 >>
rect 54 114 55 115 
<< m2c >>
rect 54 114 55 115 
<< m1 >>
rect 54 114 55 115 
<< m2 >>
rect 54 114 55 115 
<< m1 >>
rect 55 114 56 115 
<< m1 >>
rect 56 114 57 115 
<< m1 >>
rect 57 114 58 115 
<< m1 >>
rect 58 114 59 115 
<< m1 >>
rect 59 114 60 115 
<< m1 >>
rect 60 114 61 115 
<< m1 >>
rect 61 114 62 115 
<< m1 >>
rect 62 114 63 115 
<< m1 >>
rect 63 114 64 115 
<< m1 >>
rect 64 114 65 115 
<< m1 >>
rect 65 114 66 115 
<< m1 >>
rect 66 114 67 115 
<< m1 >>
rect 67 114 68 115 
<< m1 >>
rect 68 114 69 115 
<< m1 >>
rect 69 114 70 115 
<< m1 >>
rect 70 114 71 115 
<< m1 >>
rect 71 114 72 115 
<< m1 >>
rect 72 114 73 115 
<< m1 >>
rect 73 114 74 115 
<< m1 >>
rect 74 114 75 115 
<< m1 >>
rect 75 114 76 115 
<< m1 >>
rect 76 114 77 115 
<< m2 >>
rect 76 114 77 115 
<< m1 >>
rect 77 114 78 115 
<< m1 >>
rect 78 114 79 115 
<< m2 >>
rect 78 114 79 115 
<< m2c >>
rect 78 114 79 115 
<< m1 >>
rect 78 114 79 115 
<< m2 >>
rect 78 114 79 115 
<< m2 >>
rect 79 114 80 115 
<< m1 >>
rect 80 114 81 115 
<< m2 >>
rect 80 114 81 115 
<< m2 >>
rect 81 114 82 115 
<< m1 >>
rect 82 114 83 115 
<< m2 >>
rect 82 114 83 115 
<< m1 >>
rect 83 114 84 115 
<< m2 >>
rect 83 114 84 115 
<< m2c >>
rect 83 114 84 115 
<< m1 >>
rect 83 114 84 115 
<< m2 >>
rect 83 114 84 115 
<< m2 >>
rect 84 114 85 115 
<< m1 >>
rect 85 114 86 115 
<< m2 >>
rect 85 114 86 115 
<< m2 >>
rect 86 114 87 115 
<< m1 >>
rect 109 114 110 115 
<< m1 >>
rect 127 114 128 115 
<< m2 >>
rect 30 115 31 116 
<< m1 >>
rect 31 115 32 116 
<< m2 >>
rect 31 115 32 116 
<< m2 >>
rect 32 115 33 116 
<< m2 >>
rect 33 115 34 116 
<< m2 >>
rect 34 115 35 116 
<< m2 >>
rect 35 115 36 116 
<< m1 >>
rect 46 115 47 116 
<< m1 >>
rect 52 115 53 116 
<< m2 >>
rect 76 115 77 116 
<< m1 >>
rect 80 115 81 116 
<< m1 >>
rect 85 115 86 116 
<< m1 >>
rect 109 115 110 116 
<< m1 >>
rect 127 115 128 116 
<< m1 >>
rect 31 116 32 117 
<< m1 >>
rect 35 116 36 117 
<< m2 >>
rect 35 116 36 117 
<< m2c >>
rect 35 116 36 117 
<< m1 >>
rect 35 116 36 117 
<< m2 >>
rect 35 116 36 117 
<< m1 >>
rect 46 116 47 117 
<< m1 >>
rect 52 116 53 117 
<< m1 >>
rect 76 116 77 117 
<< m2 >>
rect 76 116 77 117 
<< m2c >>
rect 76 116 77 117 
<< m1 >>
rect 76 116 77 117 
<< m2 >>
rect 76 116 77 117 
<< m1 >>
rect 80 116 81 117 
<< m1 >>
rect 85 116 86 117 
<< m1 >>
rect 109 116 110 117 
<< m1 >>
rect 127 116 128 117 
<< m1 >>
rect 31 117 32 118 
<< m1 >>
rect 35 117 36 118 
<< m1 >>
rect 46 117 47 118 
<< m1 >>
rect 52 117 53 118 
<< m1 >>
rect 76 117 77 118 
<< m1 >>
rect 80 117 81 118 
<< m1 >>
rect 85 117 86 118 
<< m1 >>
rect 109 117 110 118 
<< m1 >>
rect 127 117 128 118 
<< m1 >>
rect 31 118 32 119 
<< m1 >>
rect 35 118 36 119 
<< m1 >>
rect 36 118 37 119 
<< m1 >>
rect 37 118 38 119 
<< m1 >>
rect 38 118 39 119 
<< m1 >>
rect 39 118 40 119 
<< m1 >>
rect 40 118 41 119 
<< m1 >>
rect 41 118 42 119 
<< m1 >>
rect 42 118 43 119 
<< m1 >>
rect 43 118 44 119 
<< m1 >>
rect 44 118 45 119 
<< m1 >>
rect 46 118 47 119 
<< m1 >>
rect 52 118 53 119 
<< m1 >>
rect 76 118 77 119 
<< m1 >>
rect 80 118 81 119 
<< m1 >>
rect 85 118 86 119 
<< m1 >>
rect 88 118 89 119 
<< m1 >>
rect 89 118 90 119 
<< m1 >>
rect 90 118 91 119 
<< m1 >>
rect 91 118 92 119 
<< m1 >>
rect 109 118 110 119 
<< m1 >>
rect 127 118 128 119 
<< m1 >>
rect 31 119 32 120 
<< m1 >>
rect 44 119 45 120 
<< m1 >>
rect 46 119 47 120 
<< m1 >>
rect 52 119 53 120 
<< m1 >>
rect 76 119 77 120 
<< m1 >>
rect 80 119 81 120 
<< m1 >>
rect 85 119 86 120 
<< m1 >>
rect 88 119 89 120 
<< m1 >>
rect 91 119 92 120 
<< m1 >>
rect 109 119 110 120 
<< m1 >>
rect 127 119 128 120 
<< pdiffusion >>
rect 30 120 31 121 
<< m1 >>
rect 31 120 32 121 
<< pdiffusion >>
rect 31 120 32 121 
<< pdiffusion >>
rect 32 120 33 121 
<< pdiffusion >>
rect 33 120 34 121 
<< pdiffusion >>
rect 34 120 35 121 
<< pdiffusion >>
rect 35 120 36 121 
<< m1 >>
rect 44 120 45 121 
<< m1 >>
rect 46 120 47 121 
<< pdiffusion >>
rect 48 120 49 121 
<< pdiffusion >>
rect 49 120 50 121 
<< pdiffusion >>
rect 50 120 51 121 
<< pdiffusion >>
rect 51 120 52 121 
<< m1 >>
rect 52 120 53 121 
<< pdiffusion >>
rect 52 120 53 121 
<< pdiffusion >>
rect 53 120 54 121 
<< m1 >>
rect 76 120 77 121 
<< m1 >>
rect 80 120 81 121 
<< pdiffusion >>
rect 84 120 85 121 
<< m1 >>
rect 85 120 86 121 
<< pdiffusion >>
rect 85 120 86 121 
<< pdiffusion >>
rect 86 120 87 121 
<< pdiffusion >>
rect 87 120 88 121 
<< m1 >>
rect 88 120 89 121 
<< pdiffusion >>
rect 88 120 89 121 
<< pdiffusion >>
rect 89 120 90 121 
<< m1 >>
rect 91 120 92 121 
<< pdiffusion >>
rect 102 120 103 121 
<< pdiffusion >>
rect 103 120 104 121 
<< pdiffusion >>
rect 104 120 105 121 
<< pdiffusion >>
rect 105 120 106 121 
<< pdiffusion >>
rect 106 120 107 121 
<< pdiffusion >>
rect 107 120 108 121 
<< m1 >>
rect 109 120 110 121 
<< pdiffusion >>
rect 120 120 121 121 
<< pdiffusion >>
rect 121 120 122 121 
<< pdiffusion >>
rect 122 120 123 121 
<< pdiffusion >>
rect 123 120 124 121 
<< pdiffusion >>
rect 124 120 125 121 
<< pdiffusion >>
rect 125 120 126 121 
<< m1 >>
rect 127 120 128 121 
<< pdiffusion >>
rect 30 121 31 122 
<< pdiffusion >>
rect 31 121 32 122 
<< pdiffusion >>
rect 32 121 33 122 
<< pdiffusion >>
rect 33 121 34 122 
<< pdiffusion >>
rect 34 121 35 122 
<< pdiffusion >>
rect 35 121 36 122 
<< m1 >>
rect 44 121 45 122 
<< m1 >>
rect 46 121 47 122 
<< pdiffusion >>
rect 48 121 49 122 
<< pdiffusion >>
rect 49 121 50 122 
<< pdiffusion >>
rect 50 121 51 122 
<< pdiffusion >>
rect 51 121 52 122 
<< pdiffusion >>
rect 52 121 53 122 
<< pdiffusion >>
rect 53 121 54 122 
<< m1 >>
rect 76 121 77 122 
<< m1 >>
rect 80 121 81 122 
<< pdiffusion >>
rect 84 121 85 122 
<< pdiffusion >>
rect 85 121 86 122 
<< pdiffusion >>
rect 86 121 87 122 
<< pdiffusion >>
rect 87 121 88 122 
<< pdiffusion >>
rect 88 121 89 122 
<< pdiffusion >>
rect 89 121 90 122 
<< m1 >>
rect 91 121 92 122 
<< pdiffusion >>
rect 102 121 103 122 
<< pdiffusion >>
rect 103 121 104 122 
<< pdiffusion >>
rect 104 121 105 122 
<< pdiffusion >>
rect 105 121 106 122 
<< pdiffusion >>
rect 106 121 107 122 
<< pdiffusion >>
rect 107 121 108 122 
<< m1 >>
rect 109 121 110 122 
<< pdiffusion >>
rect 120 121 121 122 
<< pdiffusion >>
rect 121 121 122 122 
<< pdiffusion >>
rect 122 121 123 122 
<< pdiffusion >>
rect 123 121 124 122 
<< pdiffusion >>
rect 124 121 125 122 
<< pdiffusion >>
rect 125 121 126 122 
<< m1 >>
rect 127 121 128 122 
<< pdiffusion >>
rect 30 122 31 123 
<< pdiffusion >>
rect 31 122 32 123 
<< pdiffusion >>
rect 32 122 33 123 
<< pdiffusion >>
rect 33 122 34 123 
<< pdiffusion >>
rect 34 122 35 123 
<< pdiffusion >>
rect 35 122 36 123 
<< m1 >>
rect 44 122 45 123 
<< m1 >>
rect 46 122 47 123 
<< pdiffusion >>
rect 48 122 49 123 
<< pdiffusion >>
rect 49 122 50 123 
<< pdiffusion >>
rect 50 122 51 123 
<< pdiffusion >>
rect 51 122 52 123 
<< pdiffusion >>
rect 52 122 53 123 
<< pdiffusion >>
rect 53 122 54 123 
<< m1 >>
rect 76 122 77 123 
<< m1 >>
rect 80 122 81 123 
<< pdiffusion >>
rect 84 122 85 123 
<< pdiffusion >>
rect 85 122 86 123 
<< pdiffusion >>
rect 86 122 87 123 
<< pdiffusion >>
rect 87 122 88 123 
<< pdiffusion >>
rect 88 122 89 123 
<< pdiffusion >>
rect 89 122 90 123 
<< m1 >>
rect 91 122 92 123 
<< pdiffusion >>
rect 102 122 103 123 
<< pdiffusion >>
rect 103 122 104 123 
<< pdiffusion >>
rect 104 122 105 123 
<< pdiffusion >>
rect 105 122 106 123 
<< pdiffusion >>
rect 106 122 107 123 
<< pdiffusion >>
rect 107 122 108 123 
<< m1 >>
rect 109 122 110 123 
<< pdiffusion >>
rect 120 122 121 123 
<< pdiffusion >>
rect 121 122 122 123 
<< pdiffusion >>
rect 122 122 123 123 
<< pdiffusion >>
rect 123 122 124 123 
<< pdiffusion >>
rect 124 122 125 123 
<< pdiffusion >>
rect 125 122 126 123 
<< m1 >>
rect 127 122 128 123 
<< pdiffusion >>
rect 30 123 31 124 
<< pdiffusion >>
rect 31 123 32 124 
<< pdiffusion >>
rect 32 123 33 124 
<< pdiffusion >>
rect 33 123 34 124 
<< pdiffusion >>
rect 34 123 35 124 
<< pdiffusion >>
rect 35 123 36 124 
<< m1 >>
rect 44 123 45 124 
<< m1 >>
rect 46 123 47 124 
<< pdiffusion >>
rect 48 123 49 124 
<< pdiffusion >>
rect 49 123 50 124 
<< pdiffusion >>
rect 50 123 51 124 
<< pdiffusion >>
rect 51 123 52 124 
<< pdiffusion >>
rect 52 123 53 124 
<< pdiffusion >>
rect 53 123 54 124 
<< m1 >>
rect 76 123 77 124 
<< m1 >>
rect 80 123 81 124 
<< pdiffusion >>
rect 84 123 85 124 
<< pdiffusion >>
rect 85 123 86 124 
<< pdiffusion >>
rect 86 123 87 124 
<< pdiffusion >>
rect 87 123 88 124 
<< pdiffusion >>
rect 88 123 89 124 
<< pdiffusion >>
rect 89 123 90 124 
<< m1 >>
rect 91 123 92 124 
<< pdiffusion >>
rect 102 123 103 124 
<< pdiffusion >>
rect 103 123 104 124 
<< pdiffusion >>
rect 104 123 105 124 
<< pdiffusion >>
rect 105 123 106 124 
<< pdiffusion >>
rect 106 123 107 124 
<< pdiffusion >>
rect 107 123 108 124 
<< m1 >>
rect 109 123 110 124 
<< pdiffusion >>
rect 120 123 121 124 
<< pdiffusion >>
rect 121 123 122 124 
<< pdiffusion >>
rect 122 123 123 124 
<< pdiffusion >>
rect 123 123 124 124 
<< pdiffusion >>
rect 124 123 125 124 
<< pdiffusion >>
rect 125 123 126 124 
<< m1 >>
rect 127 123 128 124 
<< pdiffusion >>
rect 30 124 31 125 
<< pdiffusion >>
rect 31 124 32 125 
<< pdiffusion >>
rect 32 124 33 125 
<< pdiffusion >>
rect 33 124 34 125 
<< pdiffusion >>
rect 34 124 35 125 
<< pdiffusion >>
rect 35 124 36 125 
<< m1 >>
rect 44 124 45 125 
<< m1 >>
rect 46 124 47 125 
<< pdiffusion >>
rect 48 124 49 125 
<< pdiffusion >>
rect 49 124 50 125 
<< pdiffusion >>
rect 50 124 51 125 
<< pdiffusion >>
rect 51 124 52 125 
<< pdiffusion >>
rect 52 124 53 125 
<< pdiffusion >>
rect 53 124 54 125 
<< m1 >>
rect 76 124 77 125 
<< m1 >>
rect 80 124 81 125 
<< pdiffusion >>
rect 84 124 85 125 
<< pdiffusion >>
rect 85 124 86 125 
<< pdiffusion >>
rect 86 124 87 125 
<< pdiffusion >>
rect 87 124 88 125 
<< pdiffusion >>
rect 88 124 89 125 
<< pdiffusion >>
rect 89 124 90 125 
<< m1 >>
rect 91 124 92 125 
<< pdiffusion >>
rect 102 124 103 125 
<< pdiffusion >>
rect 103 124 104 125 
<< pdiffusion >>
rect 104 124 105 125 
<< pdiffusion >>
rect 105 124 106 125 
<< pdiffusion >>
rect 106 124 107 125 
<< pdiffusion >>
rect 107 124 108 125 
<< m1 >>
rect 109 124 110 125 
<< pdiffusion >>
rect 120 124 121 125 
<< pdiffusion >>
rect 121 124 122 125 
<< pdiffusion >>
rect 122 124 123 125 
<< pdiffusion >>
rect 123 124 124 125 
<< pdiffusion >>
rect 124 124 125 125 
<< pdiffusion >>
rect 125 124 126 125 
<< m1 >>
rect 127 124 128 125 
<< pdiffusion >>
rect 30 125 31 126 
<< m1 >>
rect 31 125 32 126 
<< pdiffusion >>
rect 31 125 32 126 
<< pdiffusion >>
rect 32 125 33 126 
<< pdiffusion >>
rect 33 125 34 126 
<< pdiffusion >>
rect 34 125 35 126 
<< pdiffusion >>
rect 35 125 36 126 
<< m1 >>
rect 44 125 45 126 
<< m1 >>
rect 46 125 47 126 
<< pdiffusion >>
rect 48 125 49 126 
<< m1 >>
rect 49 125 50 126 
<< pdiffusion >>
rect 49 125 50 126 
<< pdiffusion >>
rect 50 125 51 126 
<< pdiffusion >>
rect 51 125 52 126 
<< pdiffusion >>
rect 52 125 53 126 
<< pdiffusion >>
rect 53 125 54 126 
<< m1 >>
rect 76 125 77 126 
<< m1 >>
rect 80 125 81 126 
<< pdiffusion >>
rect 84 125 85 126 
<< pdiffusion >>
rect 85 125 86 126 
<< pdiffusion >>
rect 86 125 87 126 
<< pdiffusion >>
rect 87 125 88 126 
<< pdiffusion >>
rect 88 125 89 126 
<< pdiffusion >>
rect 89 125 90 126 
<< m1 >>
rect 91 125 92 126 
<< pdiffusion >>
rect 102 125 103 126 
<< m1 >>
rect 103 125 104 126 
<< pdiffusion >>
rect 103 125 104 126 
<< pdiffusion >>
rect 104 125 105 126 
<< pdiffusion >>
rect 105 125 106 126 
<< m1 >>
rect 106 125 107 126 
<< pdiffusion >>
rect 106 125 107 126 
<< pdiffusion >>
rect 107 125 108 126 
<< m1 >>
rect 109 125 110 126 
<< pdiffusion >>
rect 120 125 121 126 
<< m1 >>
rect 121 125 122 126 
<< pdiffusion >>
rect 121 125 122 126 
<< pdiffusion >>
rect 122 125 123 126 
<< pdiffusion >>
rect 123 125 124 126 
<< pdiffusion >>
rect 124 125 125 126 
<< pdiffusion >>
rect 125 125 126 126 
<< m1 >>
rect 127 125 128 126 
<< m1 >>
rect 31 126 32 127 
<< m1 >>
rect 44 126 45 127 
<< m1 >>
rect 46 126 47 127 
<< m1 >>
rect 49 126 50 127 
<< m1 >>
rect 76 126 77 127 
<< m1 >>
rect 80 126 81 127 
<< m1 >>
rect 91 126 92 127 
<< m1 >>
rect 103 126 104 127 
<< m1 >>
rect 106 126 107 127 
<< m1 >>
rect 109 126 110 127 
<< m1 >>
rect 121 126 122 127 
<< m1 >>
rect 127 126 128 127 
<< m1 >>
rect 31 127 32 128 
<< m1 >>
rect 44 127 45 128 
<< m1 >>
rect 46 127 47 128 
<< m1 >>
rect 47 127 48 128 
<< m1 >>
rect 48 127 49 128 
<< m1 >>
rect 49 127 50 128 
<< m1 >>
rect 76 127 77 128 
<< m1 >>
rect 80 127 81 128 
<< m1 >>
rect 91 127 92 128 
<< m1 >>
rect 103 127 104 128 
<< m1 >>
rect 106 127 107 128 
<< m2 >>
rect 107 127 108 128 
<< m1 >>
rect 108 127 109 128 
<< m2 >>
rect 108 127 109 128 
<< m2c >>
rect 108 127 109 128 
<< m1 >>
rect 108 127 109 128 
<< m2 >>
rect 108 127 109 128 
<< m1 >>
rect 109 127 110 128 
<< m1 >>
rect 121 127 122 128 
<< m1 >>
rect 127 127 128 128 
<< m1 >>
rect 31 128 32 129 
<< m1 >>
rect 32 128 33 129 
<< m1 >>
rect 33 128 34 129 
<< m1 >>
rect 34 128 35 129 
<< m1 >>
rect 35 128 36 129 
<< m1 >>
rect 36 128 37 129 
<< m1 >>
rect 37 128 38 129 
<< m1 >>
rect 38 128 39 129 
<< m1 >>
rect 39 128 40 129 
<< m1 >>
rect 40 128 41 129 
<< m1 >>
rect 41 128 42 129 
<< m1 >>
rect 42 128 43 129 
<< m2 >>
rect 42 128 43 129 
<< m2c >>
rect 42 128 43 129 
<< m1 >>
rect 42 128 43 129 
<< m2 >>
rect 42 128 43 129 
<< m2 >>
rect 43 128 44 129 
<< m1 >>
rect 44 128 45 129 
<< m1 >>
rect 76 128 77 129 
<< m1 >>
rect 80 128 81 129 
<< m1 >>
rect 86 128 87 129 
<< m2 >>
rect 86 128 87 129 
<< m2c >>
rect 86 128 87 129 
<< m1 >>
rect 86 128 87 129 
<< m2 >>
rect 86 128 87 129 
<< m1 >>
rect 87 128 88 129 
<< m1 >>
rect 88 128 89 129 
<< m1 >>
rect 89 128 90 129 
<< m1 >>
rect 90 128 91 129 
<< m1 >>
rect 91 128 92 129 
<< m1 >>
rect 103 128 104 129 
<< m1 >>
rect 104 128 105 129 
<< m2 >>
rect 104 128 105 129 
<< m2c >>
rect 104 128 105 129 
<< m1 >>
rect 104 128 105 129 
<< m2 >>
rect 104 128 105 129 
<< m2 >>
rect 105 128 106 129 
<< m1 >>
rect 106 128 107 129 
<< m2 >>
rect 106 128 107 129 
<< m2 >>
rect 107 128 108 129 
<< m1 >>
rect 121 128 122 129 
<< m1 >>
rect 122 128 123 129 
<< m1 >>
rect 123 128 124 129 
<< m1 >>
rect 124 128 125 129 
<< m1 >>
rect 125 128 126 129 
<< m1 >>
rect 126 128 127 129 
<< m1 >>
rect 127 128 128 129 
<< m2 >>
rect 43 129 44 130 
<< m1 >>
rect 44 129 45 130 
<< m1 >>
rect 76 129 77 130 
<< m1 >>
rect 80 129 81 130 
<< m2 >>
rect 86 129 87 130 
<< m1 >>
rect 106 129 107 130 
<< m2 >>
rect 43 130 44 131 
<< m1 >>
rect 44 130 45 131 
<< m2 >>
rect 44 130 45 131 
<< m1 >>
rect 45 130 46 131 
<< m2 >>
rect 45 130 46 131 
<< m1 >>
rect 46 130 47 131 
<< m2 >>
rect 46 130 47 131 
<< m1 >>
rect 47 130 48 131 
<< m2 >>
rect 47 130 48 131 
<< m1 >>
rect 48 130 49 131 
<< m2 >>
rect 48 130 49 131 
<< m1 >>
rect 49 130 50 131 
<< m2 >>
rect 49 130 50 131 
<< m1 >>
rect 50 130 51 131 
<< m2 >>
rect 50 130 51 131 
<< m1 >>
rect 51 130 52 131 
<< m2 >>
rect 51 130 52 131 
<< m1 >>
rect 52 130 53 131 
<< m2 >>
rect 52 130 53 131 
<< m1 >>
rect 53 130 54 131 
<< m2 >>
rect 53 130 54 131 
<< m1 >>
rect 54 130 55 131 
<< m2 >>
rect 54 130 55 131 
<< m1 >>
rect 55 130 56 131 
<< m2 >>
rect 55 130 56 131 
<< m1 >>
rect 56 130 57 131 
<< m2 >>
rect 56 130 57 131 
<< m1 >>
rect 57 130 58 131 
<< m2 >>
rect 57 130 58 131 
<< m1 >>
rect 58 130 59 131 
<< m2 >>
rect 58 130 59 131 
<< m1 >>
rect 59 130 60 131 
<< m2 >>
rect 59 130 60 131 
<< m1 >>
rect 60 130 61 131 
<< m2 >>
rect 60 130 61 131 
<< m1 >>
rect 61 130 62 131 
<< m2 >>
rect 61 130 62 131 
<< m1 >>
rect 62 130 63 131 
<< m2 >>
rect 62 130 63 131 
<< m1 >>
rect 63 130 64 131 
<< m2 >>
rect 63 130 64 131 
<< m1 >>
rect 64 130 65 131 
<< m2 >>
rect 64 130 65 131 
<< m1 >>
rect 65 130 66 131 
<< m2 >>
rect 65 130 66 131 
<< m1 >>
rect 66 130 67 131 
<< m2 >>
rect 66 130 67 131 
<< m1 >>
rect 67 130 68 131 
<< m2 >>
rect 67 130 68 131 
<< m1 >>
rect 68 130 69 131 
<< m2 >>
rect 68 130 69 131 
<< m1 >>
rect 69 130 70 131 
<< m2 >>
rect 69 130 70 131 
<< m1 >>
rect 70 130 71 131 
<< m2 >>
rect 70 130 71 131 
<< m1 >>
rect 71 130 72 131 
<< m2 >>
rect 71 130 72 131 
<< m1 >>
rect 72 130 73 131 
<< m2 >>
rect 72 130 73 131 
<< m1 >>
rect 73 130 74 131 
<< m2 >>
rect 73 130 74 131 
<< m1 >>
rect 74 130 75 131 
<< m2 >>
rect 74 130 75 131 
<< m1 >>
rect 75 130 76 131 
<< m2 >>
rect 75 130 76 131 
<< m1 >>
rect 76 130 77 131 
<< m2 >>
rect 76 130 77 131 
<< m2 >>
rect 77 130 78 131 
<< m1 >>
rect 78 130 79 131 
<< m2 >>
rect 78 130 79 131 
<< m2c >>
rect 78 130 79 131 
<< m1 >>
rect 78 130 79 131 
<< m2 >>
rect 78 130 79 131 
<< m2 >>
rect 79 130 80 131 
<< m1 >>
rect 80 130 81 131 
<< m2 >>
rect 80 130 81 131 
<< m1 >>
rect 81 130 82 131 
<< m2 >>
rect 81 130 82 131 
<< m1 >>
rect 82 130 83 131 
<< m2 >>
rect 82 130 83 131 
<< m1 >>
rect 83 130 84 131 
<< m2 >>
rect 83 130 84 131 
<< m1 >>
rect 84 130 85 131 
<< m2 >>
rect 84 130 85 131 
<< m1 >>
rect 85 130 86 131 
<< m2 >>
rect 85 130 86 131 
<< m1 >>
rect 86 130 87 131 
<< m2 >>
rect 86 130 87 131 
<< m1 >>
rect 87 130 88 131 
<< m1 >>
rect 88 130 89 131 
<< m1 >>
rect 89 130 90 131 
<< m1 >>
rect 90 130 91 131 
<< m1 >>
rect 91 130 92 131 
<< m1 >>
rect 92 130 93 131 
<< m1 >>
rect 93 130 94 131 
<< m1 >>
rect 94 130 95 131 
<< m1 >>
rect 95 130 96 131 
<< m1 >>
rect 96 130 97 131 
<< m1 >>
rect 97 130 98 131 
<< m1 >>
rect 98 130 99 131 
<< m1 >>
rect 99 130 100 131 
<< m1 >>
rect 100 130 101 131 
<< m1 >>
rect 101 130 102 131 
<< m1 >>
rect 102 130 103 131 
<< m1 >>
rect 103 130 104 131 
<< m1 >>
rect 104 130 105 131 
<< m1 >>
rect 105 130 106 131 
<< m1 >>
rect 106 130 107 131 
<< labels >>
rlabel pdiffusion 139 84 140 85  0 t = 1
rlabel pdiffusion 142 84 143 85  0 t = 2
rlabel pdiffusion 139 89 140 90  0 t = 3
rlabel pdiffusion 142 89 143 90  0 t = 4
rlabel pdiffusion 138 84 144 90 0 cell no = 1
<< m1 >>
rect 139 84 140 85 
rect 142 84 143 85 
rect 139 89 140 90 
rect 142 89 143 90 
<< m2 >>
rect 139 84 140 85 
rect 142 84 143 85 
rect 139 89 140 90 
rect 142 89 143 90 
<< m2c >>
rect 139 84 140 85 
rect 142 84 143 85 
rect 139 89 140 90 
rect 142 89 143 90 
<< labels >>
rlabel pdiffusion 31 30 32 31  0 t = 1
rlabel pdiffusion 34 30 35 31  0 t = 2
rlabel pdiffusion 31 35 32 36  0 t = 3
rlabel pdiffusion 34 35 35 36  0 t = 4
rlabel pdiffusion 30 30 36 36 0 cell no = 2
<< m1 >>
rect 31 30 32 31 
rect 34 30 35 31 
rect 31 35 32 36 
rect 34 35 35 36 
<< m2 >>
rect 31 30 32 31 
rect 34 30 35 31 
rect 31 35 32 36 
rect 34 35 35 36 
<< m2c >>
rect 31 30 32 31 
rect 34 30 35 31 
rect 31 35 32 36 
rect 34 35 35 36 
<< labels >>
rlabel pdiffusion 49 30 50 31  0 t = 1
rlabel pdiffusion 52 30 53 31  0 t = 2
rlabel pdiffusion 49 35 50 36  0 t = 3
rlabel pdiffusion 52 35 53 36  0 t = 4
rlabel pdiffusion 48 30 54 36 0 cell no = 3
<< m1 >>
rect 49 30 50 31 
rect 52 30 53 31 
rect 49 35 50 36 
rect 52 35 53 36 
<< m2 >>
rect 49 30 50 31 
rect 52 30 53 31 
rect 49 35 50 36 
rect 52 35 53 36 
<< m2c >>
rect 49 30 50 31 
rect 52 30 53 31 
rect 49 35 50 36 
rect 52 35 53 36 
<< labels >>
rlabel pdiffusion 49 66 50 67  0 t = 1
rlabel pdiffusion 52 66 53 67  0 t = 2
rlabel pdiffusion 49 71 50 72  0 t = 3
rlabel pdiffusion 52 71 53 72  0 t = 4
rlabel pdiffusion 48 66 54 72 0 cell no = 4
<< m1 >>
rect 49 66 50 67 
rect 52 66 53 67 
rect 49 71 50 72 
rect 52 71 53 72 
<< m2 >>
rect 49 66 50 67 
rect 52 66 53 67 
rect 49 71 50 72 
rect 52 71 53 72 
<< m2c >>
rect 49 66 50 67 
rect 52 66 53 67 
rect 49 71 50 72 
rect 52 71 53 72 
<< labels >>
rlabel pdiffusion 13 102 14 103  0 t = 1
rlabel pdiffusion 16 102 17 103  0 t = 2
rlabel pdiffusion 13 107 14 108  0 t = 3
rlabel pdiffusion 16 107 17 108  0 t = 4
rlabel pdiffusion 12 102 18 108 0 cell no = 5
<< m1 >>
rect 13 102 14 103 
rect 16 102 17 103 
rect 13 107 14 108 
rect 16 107 17 108 
<< m2 >>
rect 13 102 14 103 
rect 16 102 17 103 
rect 13 107 14 108 
rect 16 107 17 108 
<< m2c >>
rect 13 102 14 103 
rect 16 102 17 103 
rect 13 107 14 108 
rect 16 107 17 108 
<< labels >>
rlabel pdiffusion 85 102 86 103  0 t = 1
rlabel pdiffusion 88 102 89 103  0 t = 2
rlabel pdiffusion 85 107 86 108  0 t = 3
rlabel pdiffusion 88 107 89 108  0 t = 4
rlabel pdiffusion 84 102 90 108 0 cell no = 6
<< m1 >>
rect 85 102 86 103 
rect 88 102 89 103 
rect 85 107 86 108 
rect 88 107 89 108 
<< m2 >>
rect 85 102 86 103 
rect 88 102 89 103 
rect 85 107 86 108 
rect 88 107 89 108 
<< m2c >>
rect 85 102 86 103 
rect 88 102 89 103 
rect 85 107 86 108 
rect 88 107 89 108 
<< labels >>
rlabel pdiffusion 103 12 104 13  0 t = 1
rlabel pdiffusion 106 12 107 13  0 t = 2
rlabel pdiffusion 103 17 104 18  0 t = 3
rlabel pdiffusion 106 17 107 18  0 t = 4
rlabel pdiffusion 102 12 108 18 0 cell no = 7
<< m1 >>
rect 103 12 104 13 
rect 106 12 107 13 
rect 103 17 104 18 
rect 106 17 107 18 
<< m2 >>
rect 103 12 104 13 
rect 106 12 107 13 
rect 103 17 104 18 
rect 106 17 107 18 
<< m2c >>
rect 103 12 104 13 
rect 106 12 107 13 
rect 103 17 104 18 
rect 106 17 107 18 
<< labels >>
rlabel pdiffusion 121 12 122 13  0 t = 1
rlabel pdiffusion 124 12 125 13  0 t = 2
rlabel pdiffusion 121 17 122 18  0 t = 3
rlabel pdiffusion 124 17 125 18  0 t = 4
rlabel pdiffusion 120 12 126 18 0 cell no = 8
<< m1 >>
rect 121 12 122 13 
rect 124 12 125 13 
rect 121 17 122 18 
rect 124 17 125 18 
<< m2 >>
rect 121 12 122 13 
rect 124 12 125 13 
rect 121 17 122 18 
rect 124 17 125 18 
<< m2c >>
rect 121 12 122 13 
rect 124 12 125 13 
rect 121 17 122 18 
rect 124 17 125 18 
<< labels >>
rlabel pdiffusion 49 12 50 13  0 t = 1
rlabel pdiffusion 52 12 53 13  0 t = 2
rlabel pdiffusion 49 17 50 18  0 t = 3
rlabel pdiffusion 52 17 53 18  0 t = 4
rlabel pdiffusion 48 12 54 18 0 cell no = 9
<< m1 >>
rect 49 12 50 13 
rect 52 12 53 13 
rect 49 17 50 18 
rect 52 17 53 18 
<< m2 >>
rect 49 12 50 13 
rect 52 12 53 13 
rect 49 17 50 18 
rect 52 17 53 18 
<< m2c >>
rect 49 12 50 13 
rect 52 12 53 13 
rect 49 17 50 18 
rect 52 17 53 18 
<< labels >>
rlabel pdiffusion 67 66 68 67  0 t = 1
rlabel pdiffusion 70 66 71 67  0 t = 2
rlabel pdiffusion 67 71 68 72  0 t = 3
rlabel pdiffusion 70 71 71 72  0 t = 4
rlabel pdiffusion 66 66 72 72 0 cell no = 10
<< m1 >>
rect 67 66 68 67 
rect 70 66 71 67 
rect 67 71 68 72 
rect 70 71 71 72 
<< m2 >>
rect 67 66 68 67 
rect 70 66 71 67 
rect 67 71 68 72 
rect 70 71 71 72 
<< m2c >>
rect 67 66 68 67 
rect 70 66 71 67 
rect 67 71 68 72 
rect 70 71 71 72 
<< labels >>
rlabel pdiffusion 121 66 122 67  0 t = 1
rlabel pdiffusion 124 66 125 67  0 t = 2
rlabel pdiffusion 121 71 122 72  0 t = 3
rlabel pdiffusion 124 71 125 72  0 t = 4
rlabel pdiffusion 120 66 126 72 0 cell no = 11
<< m1 >>
rect 121 66 122 67 
rect 124 66 125 67 
rect 121 71 122 72 
rect 124 71 125 72 
<< m2 >>
rect 121 66 122 67 
rect 124 66 125 67 
rect 121 71 122 72 
rect 124 71 125 72 
<< m2c >>
rect 121 66 122 67 
rect 124 66 125 67 
rect 121 71 122 72 
rect 124 71 125 72 
<< labels >>
rlabel pdiffusion 67 30 68 31  0 t = 1
rlabel pdiffusion 70 30 71 31  0 t = 2
rlabel pdiffusion 67 35 68 36  0 t = 3
rlabel pdiffusion 70 35 71 36  0 t = 4
rlabel pdiffusion 66 30 72 36 0 cell no = 12
<< m1 >>
rect 67 30 68 31 
rect 70 30 71 31 
rect 67 35 68 36 
rect 70 35 71 36 
<< m2 >>
rect 67 30 68 31 
rect 70 30 71 31 
rect 67 35 68 36 
rect 70 35 71 36 
<< m2c >>
rect 67 30 68 31 
rect 70 30 71 31 
rect 67 35 68 36 
rect 70 35 71 36 
<< labels >>
rlabel pdiffusion 67 48 68 49  0 t = 1
rlabel pdiffusion 70 48 71 49  0 t = 2
rlabel pdiffusion 67 53 68 54  0 t = 3
rlabel pdiffusion 70 53 71 54  0 t = 4
rlabel pdiffusion 66 48 72 54 0 cell no = 13
<< m1 >>
rect 67 48 68 49 
rect 70 48 71 49 
rect 67 53 68 54 
rect 70 53 71 54 
<< m2 >>
rect 67 48 68 49 
rect 70 48 71 49 
rect 67 53 68 54 
rect 70 53 71 54 
<< m2c >>
rect 67 48 68 49 
rect 70 48 71 49 
rect 67 53 68 54 
rect 70 53 71 54 
<< labels >>
rlabel pdiffusion 13 30 14 31  0 t = 1
rlabel pdiffusion 16 30 17 31  0 t = 2
rlabel pdiffusion 13 35 14 36  0 t = 3
rlabel pdiffusion 16 35 17 36  0 t = 4
rlabel pdiffusion 12 30 18 36 0 cell no = 14
<< m1 >>
rect 13 30 14 31 
rect 16 30 17 31 
rect 13 35 14 36 
rect 16 35 17 36 
<< m2 >>
rect 13 30 14 31 
rect 16 30 17 31 
rect 13 35 14 36 
rect 16 35 17 36 
<< m2c >>
rect 13 30 14 31 
rect 16 30 17 31 
rect 13 35 14 36 
rect 16 35 17 36 
<< labels >>
rlabel pdiffusion 103 48 104 49  0 t = 1
rlabel pdiffusion 106 48 107 49  0 t = 2
rlabel pdiffusion 103 53 104 54  0 t = 3
rlabel pdiffusion 106 53 107 54  0 t = 4
rlabel pdiffusion 102 48 108 54 0 cell no = 15
<< m1 >>
rect 103 48 104 49 
rect 106 48 107 49 
rect 103 53 104 54 
rect 106 53 107 54 
<< m2 >>
rect 103 48 104 49 
rect 106 48 107 49 
rect 103 53 104 54 
rect 106 53 107 54 
<< m2c >>
rect 103 48 104 49 
rect 106 48 107 49 
rect 103 53 104 54 
rect 106 53 107 54 
<< labels >>
rlabel pdiffusion 85 66 86 67  0 t = 1
rlabel pdiffusion 88 66 89 67  0 t = 2
rlabel pdiffusion 85 71 86 72  0 t = 3
rlabel pdiffusion 88 71 89 72  0 t = 4
rlabel pdiffusion 84 66 90 72 0 cell no = 16
<< m1 >>
rect 85 66 86 67 
rect 88 66 89 67 
rect 85 71 86 72 
rect 88 71 89 72 
<< m2 >>
rect 85 66 86 67 
rect 88 66 89 67 
rect 85 71 86 72 
rect 88 71 89 72 
<< m2c >>
rect 85 66 86 67 
rect 88 66 89 67 
rect 85 71 86 72 
rect 88 71 89 72 
<< labels >>
rlabel pdiffusion 13 66 14 67  0 t = 1
rlabel pdiffusion 16 66 17 67  0 t = 2
rlabel pdiffusion 13 71 14 72  0 t = 3
rlabel pdiffusion 16 71 17 72  0 t = 4
rlabel pdiffusion 12 66 18 72 0 cell no = 17
<< m1 >>
rect 13 66 14 67 
rect 16 66 17 67 
rect 13 71 14 72 
rect 16 71 17 72 
<< m2 >>
rect 13 66 14 67 
rect 16 66 17 67 
rect 13 71 14 72 
rect 16 71 17 72 
<< m2c >>
rect 13 66 14 67 
rect 16 66 17 67 
rect 13 71 14 72 
rect 16 71 17 72 
<< labels >>
rlabel pdiffusion 31 66 32 67  0 t = 1
rlabel pdiffusion 34 66 35 67  0 t = 2
rlabel pdiffusion 31 71 32 72  0 t = 3
rlabel pdiffusion 34 71 35 72  0 t = 4
rlabel pdiffusion 30 66 36 72 0 cell no = 18
<< m1 >>
rect 31 66 32 67 
rect 34 66 35 67 
rect 31 71 32 72 
rect 34 71 35 72 
<< m2 >>
rect 31 66 32 67 
rect 34 66 35 67 
rect 31 71 32 72 
rect 34 71 35 72 
<< m2c >>
rect 31 66 32 67 
rect 34 66 35 67 
rect 31 71 32 72 
rect 34 71 35 72 
<< labels >>
rlabel pdiffusion 13 12 14 13  0 t = 1
rlabel pdiffusion 16 12 17 13  0 t = 2
rlabel pdiffusion 13 17 14 18  0 t = 3
rlabel pdiffusion 16 17 17 18  0 t = 4
rlabel pdiffusion 12 12 18 18 0 cell no = 19
<< m1 >>
rect 13 12 14 13 
rect 16 12 17 13 
rect 13 17 14 18 
rect 16 17 17 18 
<< m2 >>
rect 13 12 14 13 
rect 16 12 17 13 
rect 13 17 14 18 
rect 16 17 17 18 
<< m2c >>
rect 13 12 14 13 
rect 16 12 17 13 
rect 13 17 14 18 
rect 16 17 17 18 
<< labels >>
rlabel pdiffusion 85 48 86 49  0 t = 1
rlabel pdiffusion 88 48 89 49  0 t = 2
rlabel pdiffusion 85 53 86 54  0 t = 3
rlabel pdiffusion 88 53 89 54  0 t = 4
rlabel pdiffusion 84 48 90 54 0 cell no = 20
<< m1 >>
rect 85 48 86 49 
rect 88 48 89 49 
rect 85 53 86 54 
rect 88 53 89 54 
<< m2 >>
rect 85 48 86 49 
rect 88 48 89 49 
rect 85 53 86 54 
rect 88 53 89 54 
<< m2c >>
rect 85 48 86 49 
rect 88 48 89 49 
rect 85 53 86 54 
rect 88 53 89 54 
<< labels >>
rlabel pdiffusion 67 102 68 103  0 t = 1
rlabel pdiffusion 70 102 71 103  0 t = 2
rlabel pdiffusion 67 107 68 108  0 t = 3
rlabel pdiffusion 70 107 71 108  0 t = 4
rlabel pdiffusion 66 102 72 108 0 cell no = 21
<< m1 >>
rect 67 102 68 103 
rect 70 102 71 103 
rect 67 107 68 108 
rect 70 107 71 108 
<< m2 >>
rect 67 102 68 103 
rect 70 102 71 103 
rect 67 107 68 108 
rect 70 107 71 108 
<< m2c >>
rect 67 102 68 103 
rect 70 102 71 103 
rect 67 107 68 108 
rect 70 107 71 108 
<< labels >>
rlabel pdiffusion 31 48 32 49  0 t = 1
rlabel pdiffusion 34 48 35 49  0 t = 2
rlabel pdiffusion 31 53 32 54  0 t = 3
rlabel pdiffusion 34 53 35 54  0 t = 4
rlabel pdiffusion 30 48 36 54 0 cell no = 22
<< m1 >>
rect 31 48 32 49 
rect 34 48 35 49 
rect 31 53 32 54 
rect 34 53 35 54 
<< m2 >>
rect 31 48 32 49 
rect 34 48 35 49 
rect 31 53 32 54 
rect 34 53 35 54 
<< m2c >>
rect 31 48 32 49 
rect 34 48 35 49 
rect 31 53 32 54 
rect 34 53 35 54 
<< labels >>
rlabel pdiffusion 139 66 140 67  0 t = 1
rlabel pdiffusion 142 66 143 67  0 t = 2
rlabel pdiffusion 139 71 140 72  0 t = 3
rlabel pdiffusion 142 71 143 72  0 t = 4
rlabel pdiffusion 138 66 144 72 0 cell no = 23
<< m1 >>
rect 139 66 140 67 
rect 142 66 143 67 
rect 139 71 140 72 
rect 142 71 143 72 
<< m2 >>
rect 139 66 140 67 
rect 142 66 143 67 
rect 139 71 140 72 
rect 142 71 143 72 
<< m2c >>
rect 139 66 140 67 
rect 142 66 143 67 
rect 139 71 140 72 
rect 142 71 143 72 
<< labels >>
rlabel pdiffusion 121 48 122 49  0 t = 1
rlabel pdiffusion 124 48 125 49  0 t = 2
rlabel pdiffusion 121 53 122 54  0 t = 3
rlabel pdiffusion 124 53 125 54  0 t = 4
rlabel pdiffusion 120 48 126 54 0 cell no = 24
<< m1 >>
rect 121 48 122 49 
rect 124 48 125 49 
rect 121 53 122 54 
rect 124 53 125 54 
<< m2 >>
rect 121 48 122 49 
rect 124 48 125 49 
rect 121 53 122 54 
rect 124 53 125 54 
<< m2c >>
rect 121 48 122 49 
rect 124 48 125 49 
rect 121 53 122 54 
rect 124 53 125 54 
<< labels >>
rlabel pdiffusion 85 12 86 13  0 t = 1
rlabel pdiffusion 88 12 89 13  0 t = 2
rlabel pdiffusion 85 17 86 18  0 t = 3
rlabel pdiffusion 88 17 89 18  0 t = 4
rlabel pdiffusion 84 12 90 18 0 cell no = 25
<< m1 >>
rect 85 12 86 13 
rect 88 12 89 13 
rect 85 17 86 18 
rect 88 17 89 18 
<< m2 >>
rect 85 12 86 13 
rect 88 12 89 13 
rect 85 17 86 18 
rect 88 17 89 18 
<< m2c >>
rect 85 12 86 13 
rect 88 12 89 13 
rect 85 17 86 18 
rect 88 17 89 18 
<< labels >>
rlabel pdiffusion 139 12 140 13  0 t = 1
rlabel pdiffusion 142 12 143 13  0 t = 2
rlabel pdiffusion 139 17 140 18  0 t = 3
rlabel pdiffusion 142 17 143 18  0 t = 4
rlabel pdiffusion 138 12 144 18 0 cell no = 26
<< m1 >>
rect 139 12 140 13 
rect 142 12 143 13 
rect 139 17 140 18 
rect 142 17 143 18 
<< m2 >>
rect 139 12 140 13 
rect 142 12 143 13 
rect 139 17 140 18 
rect 142 17 143 18 
<< m2c >>
rect 139 12 140 13 
rect 142 12 143 13 
rect 139 17 140 18 
rect 142 17 143 18 
<< labels >>
rlabel pdiffusion 121 102 122 103  0 t = 1
rlabel pdiffusion 124 102 125 103  0 t = 2
rlabel pdiffusion 121 107 122 108  0 t = 3
rlabel pdiffusion 124 107 125 108  0 t = 4
rlabel pdiffusion 120 102 126 108 0 cell no = 27
<< m1 >>
rect 121 102 122 103 
rect 124 102 125 103 
rect 121 107 122 108 
rect 124 107 125 108 
<< m2 >>
rect 121 102 122 103 
rect 124 102 125 103 
rect 121 107 122 108 
rect 124 107 125 108 
<< m2c >>
rect 121 102 122 103 
rect 124 102 125 103 
rect 121 107 122 108 
rect 124 107 125 108 
<< labels >>
rlabel pdiffusion 13 48 14 49  0 t = 1
rlabel pdiffusion 16 48 17 49  0 t = 2
rlabel pdiffusion 13 53 14 54  0 t = 3
rlabel pdiffusion 16 53 17 54  0 t = 4
rlabel pdiffusion 12 48 18 54 0 cell no = 28
<< m1 >>
rect 13 48 14 49 
rect 16 48 17 49 
rect 13 53 14 54 
rect 16 53 17 54 
<< m2 >>
rect 13 48 14 49 
rect 16 48 17 49 
rect 13 53 14 54 
rect 16 53 17 54 
<< m2c >>
rect 13 48 14 49 
rect 16 48 17 49 
rect 13 53 14 54 
rect 16 53 17 54 
<< labels >>
rlabel pdiffusion 103 30 104 31  0 t = 1
rlabel pdiffusion 106 30 107 31  0 t = 2
rlabel pdiffusion 103 35 104 36  0 t = 3
rlabel pdiffusion 106 35 107 36  0 t = 4
rlabel pdiffusion 102 30 108 36 0 cell no = 29
<< m1 >>
rect 103 30 104 31 
rect 106 30 107 31 
rect 103 35 104 36 
rect 106 35 107 36 
<< m2 >>
rect 103 30 104 31 
rect 106 30 107 31 
rect 103 35 104 36 
rect 106 35 107 36 
<< m2c >>
rect 103 30 104 31 
rect 106 30 107 31 
rect 103 35 104 36 
rect 106 35 107 36 
<< labels >>
rlabel pdiffusion 49 102 50 103  0 t = 1
rlabel pdiffusion 52 102 53 103  0 t = 2
rlabel pdiffusion 49 107 50 108  0 t = 3
rlabel pdiffusion 52 107 53 108  0 t = 4
rlabel pdiffusion 48 102 54 108 0 cell no = 30
<< m1 >>
rect 49 102 50 103 
rect 52 102 53 103 
rect 49 107 50 108 
rect 52 107 53 108 
<< m2 >>
rect 49 102 50 103 
rect 52 102 53 103 
rect 49 107 50 108 
rect 52 107 53 108 
<< m2c >>
rect 49 102 50 103 
rect 52 102 53 103 
rect 49 107 50 108 
rect 52 107 53 108 
<< labels >>
rlabel pdiffusion 121 30 122 31  0 t = 1
rlabel pdiffusion 124 30 125 31  0 t = 2
rlabel pdiffusion 121 35 122 36  0 t = 3
rlabel pdiffusion 124 35 125 36  0 t = 4
rlabel pdiffusion 120 30 126 36 0 cell no = 31
<< m1 >>
rect 121 30 122 31 
rect 124 30 125 31 
rect 121 35 122 36 
rect 124 35 125 36 
<< m2 >>
rect 121 30 122 31 
rect 124 30 125 31 
rect 121 35 122 36 
rect 124 35 125 36 
<< m2c >>
rect 121 30 122 31 
rect 124 30 125 31 
rect 121 35 122 36 
rect 124 35 125 36 
<< labels >>
rlabel pdiffusion 103 84 104 85  0 t = 1
rlabel pdiffusion 106 84 107 85  0 t = 2
rlabel pdiffusion 103 89 104 90  0 t = 3
rlabel pdiffusion 106 89 107 90  0 t = 4
rlabel pdiffusion 102 84 108 90 0 cell no = 32
<< m1 >>
rect 103 84 104 85 
rect 106 84 107 85 
rect 103 89 104 90 
rect 106 89 107 90 
<< m2 >>
rect 103 84 104 85 
rect 106 84 107 85 
rect 103 89 104 90 
rect 106 89 107 90 
<< m2c >>
rect 103 84 104 85 
rect 106 84 107 85 
rect 103 89 104 90 
rect 106 89 107 90 
<< labels >>
rlabel pdiffusion 49 48 50 49  0 t = 1
rlabel pdiffusion 52 48 53 49  0 t = 2
rlabel pdiffusion 49 53 50 54  0 t = 3
rlabel pdiffusion 52 53 53 54  0 t = 4
rlabel pdiffusion 48 48 54 54 0 cell no = 33
<< m1 >>
rect 49 48 50 49 
rect 52 48 53 49 
rect 49 53 50 54 
rect 52 53 53 54 
<< m2 >>
rect 49 48 50 49 
rect 52 48 53 49 
rect 49 53 50 54 
rect 52 53 53 54 
<< m2c >>
rect 49 48 50 49 
rect 52 48 53 49 
rect 49 53 50 54 
rect 52 53 53 54 
<< labels >>
rlabel pdiffusion 103 102 104 103  0 t = 1
rlabel pdiffusion 106 102 107 103  0 t = 2
rlabel pdiffusion 103 107 104 108  0 t = 3
rlabel pdiffusion 106 107 107 108  0 t = 4
rlabel pdiffusion 102 102 108 108 0 cell no = 34
<< m1 >>
rect 103 102 104 103 
rect 106 102 107 103 
rect 103 107 104 108 
rect 106 107 107 108 
<< m2 >>
rect 103 102 104 103 
rect 106 102 107 103 
rect 103 107 104 108 
rect 106 107 107 108 
<< m2c >>
rect 103 102 104 103 
rect 106 102 107 103 
rect 103 107 104 108 
rect 106 107 107 108 
<< labels >>
rlabel pdiffusion 31 102 32 103  0 t = 1
rlabel pdiffusion 34 102 35 103  0 t = 2
rlabel pdiffusion 31 107 32 108  0 t = 3
rlabel pdiffusion 34 107 35 108  0 t = 4
rlabel pdiffusion 30 102 36 108 0 cell no = 35
<< m1 >>
rect 31 102 32 103 
rect 34 102 35 103 
rect 31 107 32 108 
rect 34 107 35 108 
<< m2 >>
rect 31 102 32 103 
rect 34 102 35 103 
rect 31 107 32 108 
rect 34 107 35 108 
<< m2c >>
rect 31 102 32 103 
rect 34 102 35 103 
rect 31 107 32 108 
rect 34 107 35 108 
<< labels >>
rlabel pdiffusion 103 66 104 67  0 t = 1
rlabel pdiffusion 106 66 107 67  0 t = 2
rlabel pdiffusion 103 71 104 72  0 t = 3
rlabel pdiffusion 106 71 107 72  0 t = 4
rlabel pdiffusion 102 66 108 72 0 cell no = 36
<< m1 >>
rect 103 66 104 67 
rect 106 66 107 67 
rect 103 71 104 72 
rect 106 71 107 72 
<< m2 >>
rect 103 66 104 67 
rect 106 66 107 67 
rect 103 71 104 72 
rect 106 71 107 72 
<< m2c >>
rect 103 66 104 67 
rect 106 66 107 67 
rect 103 71 104 72 
rect 106 71 107 72 
<< labels >>
rlabel pdiffusion 49 120 50 121  0 t = 1
rlabel pdiffusion 52 120 53 121  0 t = 2
rlabel pdiffusion 49 125 50 126  0 t = 3
rlabel pdiffusion 52 125 53 126  0 t = 4
rlabel pdiffusion 48 120 54 126 0 cell no = 37
<< m1 >>
rect 49 120 50 121 
rect 52 120 53 121 
rect 49 125 50 126 
rect 52 125 53 126 
<< m2 >>
rect 49 120 50 121 
rect 52 120 53 121 
rect 49 125 50 126 
rect 52 125 53 126 
<< m2c >>
rect 49 120 50 121 
rect 52 120 53 121 
rect 49 125 50 126 
rect 52 125 53 126 
<< labels >>
rlabel pdiffusion 49 84 50 85  0 t = 1
rlabel pdiffusion 52 84 53 85  0 t = 2
rlabel pdiffusion 49 89 50 90  0 t = 3
rlabel pdiffusion 52 89 53 90  0 t = 4
rlabel pdiffusion 48 84 54 90 0 cell no = 38
<< m1 >>
rect 49 84 50 85 
rect 52 84 53 85 
rect 49 89 50 90 
rect 52 89 53 90 
<< m2 >>
rect 49 84 50 85 
rect 52 84 53 85 
rect 49 89 50 90 
rect 52 89 53 90 
<< m2c >>
rect 49 84 50 85 
rect 52 84 53 85 
rect 49 89 50 90 
rect 52 89 53 90 
<< labels >>
rlabel pdiffusion 139 48 140 49  0 t = 1
rlabel pdiffusion 142 48 143 49  0 t = 2
rlabel pdiffusion 139 53 140 54  0 t = 3
rlabel pdiffusion 142 53 143 54  0 t = 4
rlabel pdiffusion 138 48 144 54 0 cell no = 39
<< m1 >>
rect 139 48 140 49 
rect 142 48 143 49 
rect 139 53 140 54 
rect 142 53 143 54 
<< m2 >>
rect 139 48 140 49 
rect 142 48 143 49 
rect 139 53 140 54 
rect 142 53 143 54 
<< m2c >>
rect 139 48 140 49 
rect 142 48 143 49 
rect 139 53 140 54 
rect 142 53 143 54 
<< labels >>
rlabel pdiffusion 31 120 32 121  0 t = 1
rlabel pdiffusion 34 120 35 121  0 t = 2
rlabel pdiffusion 31 125 32 126  0 t = 3
rlabel pdiffusion 34 125 35 126  0 t = 4
rlabel pdiffusion 30 120 36 126 0 cell no = 40
<< m1 >>
rect 31 120 32 121 
rect 34 120 35 121 
rect 31 125 32 126 
rect 34 125 35 126 
<< m2 >>
rect 31 120 32 121 
rect 34 120 35 121 
rect 31 125 32 126 
rect 34 125 35 126 
<< m2c >>
rect 31 120 32 121 
rect 34 120 35 121 
rect 31 125 32 126 
rect 34 125 35 126 
<< labels >>
rlabel pdiffusion 85 120 86 121  0 t = 1
rlabel pdiffusion 88 120 89 121  0 t = 2
rlabel pdiffusion 85 125 86 126  0 t = 3
rlabel pdiffusion 88 125 89 126  0 t = 4
rlabel pdiffusion 84 120 90 126 0 cell no = 41
<< m1 >>
rect 85 120 86 121 
rect 88 120 89 121 
rect 85 125 86 126 
rect 88 125 89 126 
<< m2 >>
rect 85 120 86 121 
rect 88 120 89 121 
rect 85 125 86 126 
rect 88 125 89 126 
<< m2c >>
rect 85 120 86 121 
rect 88 120 89 121 
rect 85 125 86 126 
rect 88 125 89 126 
<< labels >>
rlabel pdiffusion 85 84 86 85  0 t = 1
rlabel pdiffusion 88 84 89 85  0 t = 2
rlabel pdiffusion 85 89 86 90  0 t = 3
rlabel pdiffusion 88 89 89 90  0 t = 4
rlabel pdiffusion 84 84 90 90 0 cell no = 42
<< m1 >>
rect 85 84 86 85 
rect 88 84 89 85 
rect 85 89 86 90 
rect 88 89 89 90 
<< m2 >>
rect 85 84 86 85 
rect 88 84 89 85 
rect 85 89 86 90 
rect 88 89 89 90 
<< m2c >>
rect 85 84 86 85 
rect 88 84 89 85 
rect 85 89 86 90 
rect 88 89 89 90 
<< labels >>
rlabel pdiffusion 103 120 104 121  0 t = 1
rlabel pdiffusion 106 120 107 121  0 t = 2
rlabel pdiffusion 103 125 104 126  0 t = 3
rlabel pdiffusion 106 125 107 126  0 t = 4
rlabel pdiffusion 102 120 108 126 0 cell no = 43
<< m1 >>
rect 103 120 104 121 
rect 106 120 107 121 
rect 103 125 104 126 
rect 106 125 107 126 
<< m2 >>
rect 103 120 104 121 
rect 106 120 107 121 
rect 103 125 104 126 
rect 106 125 107 126 
<< m2c >>
rect 103 120 104 121 
rect 106 120 107 121 
rect 103 125 104 126 
rect 106 125 107 126 
<< labels >>
rlabel pdiffusion 67 84 68 85  0 t = 1
rlabel pdiffusion 70 84 71 85  0 t = 2
rlabel pdiffusion 67 89 68 90  0 t = 3
rlabel pdiffusion 70 89 71 90  0 t = 4
rlabel pdiffusion 66 84 72 90 0 cell no = 44
<< m1 >>
rect 67 84 68 85 
rect 70 84 71 85 
rect 67 89 68 90 
rect 70 89 71 90 
<< m2 >>
rect 67 84 68 85 
rect 70 84 71 85 
rect 67 89 68 90 
rect 70 89 71 90 
<< m2c >>
rect 67 84 68 85 
rect 70 84 71 85 
rect 67 89 68 90 
rect 70 89 71 90 
<< labels >>
rlabel pdiffusion 13 84 14 85  0 t = 1
rlabel pdiffusion 16 84 17 85  0 t = 2
rlabel pdiffusion 13 89 14 90  0 t = 3
rlabel pdiffusion 16 89 17 90  0 t = 4
rlabel pdiffusion 12 84 18 90 0 cell no = 45
<< m1 >>
rect 13 84 14 85 
rect 16 84 17 85 
rect 13 89 14 90 
rect 16 89 17 90 
<< m2 >>
rect 13 84 14 85 
rect 16 84 17 85 
rect 13 89 14 90 
rect 16 89 17 90 
<< m2c >>
rect 13 84 14 85 
rect 16 84 17 85 
rect 13 89 14 90 
rect 16 89 17 90 
<< labels >>
rlabel pdiffusion 67 12 68 13  0 t = 1
rlabel pdiffusion 70 12 71 13  0 t = 2
rlabel pdiffusion 67 17 68 18  0 t = 3
rlabel pdiffusion 70 17 71 18  0 t = 4
rlabel pdiffusion 66 12 72 18 0 cell no = 46
<< m1 >>
rect 67 12 68 13 
rect 70 12 71 13 
rect 67 17 68 18 
rect 70 17 71 18 
<< m2 >>
rect 67 12 68 13 
rect 70 12 71 13 
rect 67 17 68 18 
rect 70 17 71 18 
<< m2c >>
rect 67 12 68 13 
rect 70 12 71 13 
rect 67 17 68 18 
rect 70 17 71 18 
<< labels >>
rlabel pdiffusion 85 30 86 31  0 t = 1
rlabel pdiffusion 88 30 89 31  0 t = 2
rlabel pdiffusion 85 35 86 36  0 t = 3
rlabel pdiffusion 88 35 89 36  0 t = 4
rlabel pdiffusion 84 30 90 36 0 cell no = 47
<< m1 >>
rect 85 30 86 31 
rect 88 30 89 31 
rect 85 35 86 36 
rect 88 35 89 36 
<< m2 >>
rect 85 30 86 31 
rect 88 30 89 31 
rect 85 35 86 36 
rect 88 35 89 36 
<< m2c >>
rect 85 30 86 31 
rect 88 30 89 31 
rect 85 35 86 36 
rect 88 35 89 36 
<< labels >>
rlabel pdiffusion 121 120 122 121  0 t = 1
rlabel pdiffusion 124 120 125 121  0 t = 2
rlabel pdiffusion 121 125 122 126  0 t = 3
rlabel pdiffusion 124 125 125 126  0 t = 4
rlabel pdiffusion 120 120 126 126 0 cell no = 48
<< m1 >>
rect 121 120 122 121 
rect 124 120 125 121 
rect 121 125 122 126 
rect 124 125 125 126 
<< m2 >>
rect 121 120 122 121 
rect 124 120 125 121 
rect 121 125 122 126 
rect 124 125 125 126 
<< m2c >>
rect 121 120 122 121 
rect 124 120 125 121 
rect 121 125 122 126 
rect 124 125 125 126 
<< labels >>
rlabel pdiffusion 139 102 140 103  0 t = 1
rlabel pdiffusion 142 102 143 103  0 t = 2
rlabel pdiffusion 139 107 140 108  0 t = 3
rlabel pdiffusion 142 107 143 108  0 t = 4
rlabel pdiffusion 138 102 144 108 0 cell no = 49
<< m1 >>
rect 139 102 140 103 
rect 142 102 143 103 
rect 139 107 140 108 
rect 142 107 143 108 
<< m2 >>
rect 139 102 140 103 
rect 142 102 143 103 
rect 139 107 140 108 
rect 142 107 143 108 
<< m2c >>
rect 139 102 140 103 
rect 142 102 143 103 
rect 139 107 140 108 
rect 142 107 143 108 
<< labels >>
rlabel pdiffusion 31 84 32 85  0 t = 1
rlabel pdiffusion 34 84 35 85  0 t = 2
rlabel pdiffusion 31 89 32 90  0 t = 3
rlabel pdiffusion 34 89 35 90  0 t = 4
rlabel pdiffusion 30 84 36 90 0 cell no = 50
<< m1 >>
rect 31 84 32 85 
rect 34 84 35 85 
rect 31 89 32 90 
rect 34 89 35 90 
<< m2 >>
rect 31 84 32 85 
rect 34 84 35 85 
rect 31 89 32 90 
rect 34 89 35 90 
<< m2c >>
rect 31 84 32 85 
rect 34 84 35 85 
rect 31 89 32 90 
rect 34 89 35 90 
<< end >> 
